------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    2020-07-16
-- Module Name:    GEM_LOADER
-- Description:    This module implements the so called gemloader module which stores the frontend firmware, and streams it to the gem logic on request.
--                 This version uses the FPGA BRAM for storing the bitfile  
------------------------------------------------------------------------------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library xpm;
use xpm.vcomponents.all;

use work.ttc_pkg.all;
use work.common_pkg.all;
use work.gem_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity promless is
    generic(
        g_MAX_SIZE_BYTES    : integer; -- NOTE: must be a multiple of 32KB (kilobytes) if g_MEMORY_PRIMITIVE is set to "ultra" (using UltraRAM)
        g_MEMORY_PRIMITIVE  : string := "ultra"
    );
    port (
        reset_i             : in  std_logic;
        
        to_gem_loader_i     : in  t_to_gem_loader;
        from_gem_loader_o   : out t_from_gem_loader;        
        
        -- IPbus
        ipb_reset_i         : in  std_logic;
        ipb_clk_i           : in  std_logic;
        ipb_miso_o          : out ipb_rbus;
        ipb_mosi_i          : in  ipb_wbus                
    );
end promless;

architecture promless_arch of promless is

    ----==== RAM signals ====----
    
    -- port A is used by the IPbus slave (write and read), and port B is used by the loader (read-only)
    
    constant RAM_ADDR_WIDTH_A : integer := 22;
    constant RAM_ADDR_WIDTH_B : integer := 24;
    
    -- Common RAM port A signals 
    signal rama_addr                : std_logic_vector(RAM_ADDR_WIDTH_A - 1 downto 0) := (others => '0');
    signal rama_din                 : std_logic_vector(31 downto 0) := (others => '0');
    signal rama_we                  : std_logic  := '0';
    signal rama_dout                : std_logic_vector(31 downto 0);

    signal rama_write_req           : std_logic;
    signal rama_read_req            : std_logic;
    signal rama_read_ready          : std_logic;
    signal rama_read_ready_pipe     : std_logic_vector(1 downto 0) := (others => '0');
    signal rama_write_addr          : std_logic_vector(RAM_ADDR_WIDTH_A - 1 downto 0) := (others => '0');
    signal rama_read_addr           : std_logic_vector(RAM_ADDR_WIDTH_A - 1 downto 0) := (others => '0');
    signal rama_reset_addr          : std_logic;

    -- port B signals
    signal ramb_addr                : std_logic_vector(RAM_ADDR_WIDTH_B - 1 downto 0) := (others => '0');
    signal ramb_dout                : std_logic_vector(7 downto 0);
    
    ----==== Loader signals ====----
    signal firmware_size            : std_logic_vector(RAM_ADDR_WIDTH_B - 1 downto 0) := (others => '0');
    signal loader_clk               : std_logic;
    signal loader_en_req            : std_logic;
    signal from_gem_loader          : t_from_gem_loader;
    signal loader_valid_pipe        : std_logic_vector(1 downto 0) := (others => '0');

    ------ Register signals begin (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    ------ Register signals end ----------------------------------------------
        
begin

    loader_clk <= to_gem_loader_i.clk;
    loader_en_req <= to_gem_loader_i.en;

    ----==== RAM instantiation ====----    

    i_gbtx_config_ram : xpm_memory_tdpram
        generic map(
            MEMORY_SIZE        => g_MAX_SIZE_BYTES,
            MEMORY_PRIMITIVE   => g_MEMORY_PRIMITIVE,
            CLOCKING_MODE      => "common_clock",
            ECC_MODE           => "no_ecc",
            MEMORY_INIT_FILE   => "none",
            MEMORY_INIT_PARAM  => "0",
            USE_MEM_INIT       => 0,
            WAKEUP_TIME        => "disable_sleep",
            AUTO_SLEEP_TIME    => 0,
            MESSAGE_CONTROL    => 0,
            WRITE_DATA_WIDTH_A => 32,
            READ_DATA_WIDTH_A  => 32,
            BYTE_WRITE_WIDTH_A => 32,
            ADDR_WIDTH_A       => RAM_ADDR_WIDTH_A,
            READ_RESET_VALUE_A => "0",
            READ_LATENCY_A     => 2,
            WRITE_MODE_A       => "no_change",
            WRITE_DATA_WIDTH_B => 8,
            READ_DATA_WIDTH_B  => 8,
            BYTE_WRITE_WIDTH_B => 8,
            ADDR_WIDTH_B       => RAM_ADDR_WIDTH_B,
            READ_RESET_VALUE_B => "0",
            READ_LATENCY_B     => 2,
            WRITE_MODE_B       => "no_change"
        )
        port map(
            sleep          => '0',
            clka           => loader_clk,
            rsta           => '0',
            ena            => '1',
            regcea         => '1',
            wea            => (others => rama_we),
            addra          => rama_addr,
            dina           => rama_din,
            injectsbiterra => '0',
            injectdbiterra => '0',
            douta          => rama_dout,
            sbiterra       => open,
            dbiterra       => open,
            clkb           => loader_clk,
            rstb           => '0',
            enb            => '1',
            regceb         => '1',
            web            => (others => '0'),
            addrb          => ramb_addr,
            dinb           => (others => '0'),
            injectsbiterrb => '0',
            injectdbiterrb => '0',
            doutb          => ramb_dout,
            sbiterrb       => open,
            dbiterrb       => open
        );

    ----==== BRAM reading / writing ====----    
    
    -- rama_din and rama_dout are connected to WRITE_DATA and READ_DATA registers
    -- whenever a write request to WRITE_DATA is done, WE is asserted and the write address is then incremented by 1
    -- same happens with the read requests
    process (loader_clk)
    begin
        if rising_edge(loader_clk) then
            if (reset_i = '1' or rama_reset_addr = '1') then
                rama_write_addr <= (others => '0');
                rama_read_addr <= (others => '0');
            else
                rama_we <= rama_write_req; 
                if (rama_write_req = '1') then
                    rama_addr <= rama_write_addr;
                end if;
                if (rama_we = '1') then
                    rama_write_addr <= std_logic_vector(unsigned(rama_write_addr) + 1);
                end if;
                
                if (rama_read_req = '1') then
                    rama_addr <= rama_read_addr;
                end if;
                if (rama_read_ready = '1') then
                    rama_read_addr <= std_logic_vector(unsigned(rama_read_addr) + 1);
                end if;
                rama_read_ready_pipe(1) <= rama_read_req;
                rama_read_ready_pipe(0) <= rama_read_ready_pipe(1);
                rama_read_ready <= rama_read_ready_pipe(0);
                
            end if;
        end if;
    end process;

    ----==== Loader ====----    

    from_gem_loader.first <= '0';
    from_gem_loader.last <= '0';
    from_gem_loader.error <= '0';

    process(loader_clk)
    begin
        if rising_edge(loader_clk) then
            if (reset_i = '1') then
                ramb_addr <= (others => '0');
                from_gem_loader.ready <= '0';
                from_gem_loader.valid <= '0';
                from_gem_loader.data <= (others => '0');
                loader_valid_pipe <= (others => '0');
            else
                
                loader_valid_pipe(0) <= loader_valid_pipe(1);
                from_gem_loader.valid <= loader_valid_pipe(0);
                from_gem_loader.data <= ramb_dout;
                
                -- IDLE
                if (ramb_addr = std_logic_vector(to_unsigned(0, RAM_ADDR_WIDTH_B))) then
                    -- request
                    if (loader_en_req = '1') then
                        loader_valid_pipe(1) <= '1';
                        ramb_addr <= std_logic_vector(unsigned(ramb_addr) + 1);
                        from_gem_loader.ready <= '0';
                    --idle
                    else
                        loader_valid_pipe(1) <= '0';
                        ramb_addr <= (others => '0');
                        from_gem_loader.ready <= '1';
                    end if;
                    
                -- DONE
                elsif (ramb_addr = firmware_size) then
                    loader_valid_pipe(1) <= '0';
                    ramb_addr <= (others => '0');
                    from_gem_loader.ready <= '1';                    
                
                -- RUNNING
                else
                    loader_valid_pipe(1) <= '1';
                    ramb_addr <= std_logic_vector(unsigned(ramb_addr) + 1);
                    from_gem_loader.ready <= '0';
                end if;
            end if;
        end if;
    end process;
        
    -- register the output
    process(loader_clk)
    begin
        if rising_edge(loader_clk) then
            from_gem_loader_o <= from_gem_loader;
        end if;
    end process;


    --===============================================================================================
    -- this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    --==== Registers end ============================================================================
    
end promless_arch;
