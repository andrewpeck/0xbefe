----------------------------------------------------------------------------------
-- Company: TAMU, a lot of this is taken from WU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date: 14.03.2023
-- Module Name: TTC_LINK_GBTX
-- Project Name:
-- Description: A special TTC receiver that can be used in labs -- it can receive a TTC stream from a standard GE2/1 GBT0 link
--              so e.g. you can have a CTP7 running GE2/1 firmware, and connect any of its OH# GBT0 link to this receiver, and the CTP7 TTC commands will be received here     
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

library UNISIM;
use UNISIM.VComponents.all;

--use work.ctp7_utils_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.common_pkg.all;
use work.ipb_addr_decode.all;
use work.registers.all;

--============================================================================
--                                                          Entity declaration
--============================================================================

entity ttc_link_gbtx is
    generic(
        g_IPB_CLK_PERIOD_NS  : integer
    );
    port(
        -- reset
        reset_i             : in  std_logic;

        -- TTC clocks
        ttc_clks_i          : in  t_ttc_clks;

        -- GBT link
        gt_gbt_rx_data_i    : in  std_logic_vector(39 downto 0);
        gt_gbt_rx_clk_i     : in  std_logic;
        gt_gbt_status_i     : in  t_mgt_status;
        gt_gbt_ctrl_o       : out t_mgt_ctrl;

        -- TTC commands
        ttc_cmds_o          : out t_ttc_cmds;
    
        -- IPbus
        ipb_reset_i         : in  std_logic;
        ipb_clk_i           : in  std_logic;
        ipb_mosi_i          : in  ipb_wbus;
        ipb_miso_o          : out ipb_rbus
    );

end ttc_link_gbtx;

--============================================================================
--                                                        Architecture section
--============================================================================
architecture behavioral of ttc_link_gbtx is

    --============================================================================
    --                                                         Signal declarations
    --============================================================================

    signal reset                    : std_logic;
    signal ext_reset_sync           : std_logic;
    signal reset_local              : std_logic;
    signal cnt_reset                : std_logic;

    signal gbt_rx_phase             : std_logic_vector(5 downto 0);
    signal gbt_rx_phase_auto        : std_logic;
    signal gbt_rx_data              : std_logic_vector(83 downto 0);
    signal gbt_status               : t_gbt_link_status;

    ------ Register signals begin (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    ------ Register signals end ----------------------------------------------
    
--============================================================================
--                                                          Architecture begin
--============================================================================

begin

    ------------- Wiring and resets -------------

    i_reset_sync: 
    entity work.synch
        generic map(
            N_STAGES => 3
        )
        port map(
            async_i => reset_i,
            clk_i   => ttc_clks_i.clk_40,
            sync_o  => ext_reset_sync
        );

    reset <= ext_reset_sync or reset_local;

    ------------- GBTX link -------------
    
    i_gbt : entity work.gbt
        generic map(
            NUM_LINKS           => 1,
            TX_OPTIMIZATION     => 0,
            RX_OPTIMIZATION     => 0, -- TODO: must be 1
            TX_ENCODING         => 0,
            RX_ENCODING_EVEN    => 0,
            RX_ENCODING_ODD     => 0,
            g_USE_RX_SYNC_FIFOS => false
        )
        port map(
            reset_i                     => reset,
            cnt_reset_i                 => cnt_reset,

            tx_frame_clk_i              => ttc_clks_i.clk_40,
            rx_frame_clk_i              => ttc_clks_i.clk_40,
            rx_word_common_clk_i        => ttc_clks_i.clk_120,
            tx_word_clk_arr_i           => (others => ttc_clks_i.clk_120),
            rx_word_clk_arr_i           => (others => gt_gbt_rx_clk_i),

            tx_we_arr_i                 => (others => '1'),
            tx_data_arr_i               => (others => (others => '0')),
            tx_bitslip_cnt_i            => (others => (others => '0')),

            rx_bitslip_cnt_i            => (others => (others => '0')),
            rx_bitslip_auto_i           => (others => '0'),
            rx_data_valid_arr_o         => open,
            rx_data_arr_o(0)            => gbt_rx_data,
            rx_data_widebus_arr_o       => open,

            mgt_status_arr_i            => (others => gt_gbt_status_i),
            mgt_ctrl_arr_o(0)           => gt_gbt_ctrl_o,
            mgt_tx_data_arr_o           => open,
            mgt_rx_data_arr_i           => (others => gt_gbt_rx_data_i),

            prbs_mode_en_i              => '0',
            link_status_arr_o(0)        => gbt_status
        );

    ------------- GBTX link -------------

    process(ttc_clks_i.clk_40)
    begin
        if rising_edge(ttc_clks_i.clk_40) then
            if reset = '1' or gbt_status.gbt_rx_ready = '0' then
                ttc_cmds_o <= TTC_CMDS_NULL;
            else
                ttc_cmds_o.l1a <= gbt_rx_data(71);
                ttc_cmds_o.bc0 <= gbt_rx_data(70);
                ttc_cmds_o.ec0 <= gbt_rx_data(69);
                ttc_cmds_o.oc0 <= gbt_rx_data(68);
                ttc_cmds_o.resync <= gbt_rx_data(67);
                ttc_cmds_o.hard_reset <= gbt_rx_data(66);
                ttc_cmds_o.calpulse <= gbt_rx_data(65);
                ttc_cmds_o.test_sync <= gbt_rx_data(64);
            end if;
        end if;
    end process;
            
    --===============================================================================================
    -- this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    --==== Registers end ==================================================ttc_receiver_gbtx===================

end behavioral;
--============================================================================
--                                                            Architecture end
--============================================================================
