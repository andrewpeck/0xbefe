------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    12:22 2016-05-10
-- Module Name:    trigger
-- Description:    This module handles everything related to sbit cluster data (link synchronization, monitoring, local triggering, matching to L1A and reporting data to DAQ)  
------------------------------------------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

library xpm;
use xpm.vcomponents.all;

use work.common_pkg.all;
use work.gem_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity oh_link_regs is
    generic(
        g_GEM_STATION       : integer;
        g_NUM_OF_OHs        : integer;
        g_NUM_GBTS_PER_OH   : integer;
        g_IPB_CLK_PERIOD_NS : integer
    );
    port(
        -- reset
        reset_i                     : in  std_logic;
        clk_i                       : in  std_logic;

        -- Link statuses
        gbt_link_status_arr_i       : in t_gbt_link_status_arr(g_NUM_OF_OHs * g_NUM_GBTS_PER_OH - 1 downto 0);
        vfat3_link_status_arr_i     : in t_oh_vfat_link_status_arr(g_NUM_OF_OHs - 1 downto 0);

        -- Control
        vfat_mask_arr_o             : out t_std24_array(g_NUM_OF_OHs - 1 downto 0);
        gbt_tx_bitslip_arr_o        : out t_std7_array(g_NUM_OF_OHs * g_NUM_GBTS_PER_OH - 1 downto 0);
        gbt_rx_bitslip_arr_o        : out t_std6_array(g_NUM_OF_OHs * g_NUM_GBTS_PER_OH - 1 downto 0);        
        gbt_rx_bitslip_auto_arr_o   : out std_logic_vector(g_NUM_OF_OHs * g_NUM_GBTS_PER_OH - 1 downto 0);        

        -- Spy link
        spy_rx_usrclk_i             : in  std_logic;
        spy_rx_data_i               : in  t_mgt_64b_rx_data;
        spy_status_i                : in  t_mgt_status;
                                    
        -- IPbus                    
        ipb_reset_i                 : in  std_logic;
        ipb_clk_i                   : in  std_logic;
        ipb_miso_o                  : out ipb_rbus;
        ipb_mosi_i                  : in  ipb_wbus
    );
end oh_link_regs;

architecture oh_link_regs_arch of oh_link_regs is
    
    signal vfat_mask_arr            : t_std24_array(g_NUM_OF_OHs - 1 downto 0);
    signal gbt_tx_bitslip_arr       : t_std7_array(g_NUM_OF_OHs * g_NUM_GBTS_PER_OH - 1 downto 0);
    signal gbt_rx_bitslip_arr       : t_std6_array(g_NUM_OF_OHs * g_NUM_GBTS_PER_OH - 1 downto 0);
    signal gbt_rx_bitslip_auto_arr  : std_logic_vector(g_NUM_OF_OHs * g_NUM_GBTS_PER_OH - 1 downto 0);
    
    signal spy_mgt_buf_ovf          : std_logic_vector(15 downto 0);
    signal spy_mgt_buf_unf          : std_logic_vector(15 downto 0);
    signal spy_not_in_table         : std_logic_vector(15 downto 0);
    signal spy_disperr              : std_logic_vector(15 downto 0);
    signal spy_clk_corr_add         : std_logic_vector(15 downto 0);
    signal spy_clk_corr_drop        : std_logic_vector(15 downto 0);

    signal spy_mgt_buf_ovf_sync     : std_logic_vector(15 downto 0);
    signal spy_mgt_buf_unf_sync     : std_logic_vector(15 downto 0);
    signal spy_not_in_table_sync    : std_logic_vector(15 downto 0);
    signal spy_disperr_sync         : std_logic_vector(15 downto 0);
    signal spy_clk_corr_add_sync    : std_logic_vector(15 downto 0);
    signal spy_clk_corr_drop_sync   : std_logic_vector(15 downto 0);
    
    ------ Register signals begin ge11 (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    ------ Register signals end ge11 ----------------------------------------------

    ------ Register signals begin ge21 (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    ------ Register signals end ge21 ----------------------------------------------

    ------ Register signals begin me0 (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    ------ Register signals end me0 ----------------------------------------------
    
begin
    
    vfat_mask_arr_o <= vfat_mask_arr;
    gbt_tx_bitslip_arr_o <= gbt_tx_bitslip_arr;
    gbt_rx_bitslip_arr_o <= gbt_rx_bitslip_arr;
    gbt_rx_bitslip_auto_arr_o <= gbt_rx_bitslip_auto_arr;
    
    --================================--
    -- Spy link counters  
    --================================--

    -- elastic buffer overflow counter
    i_cnt_spy_mgt_buf_ovf : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => spy_rx_usrclk_i,
            reset_i   => reset_i,
            en_i      => (spy_status_i.rxbufstatus(2)) and (spy_status_i.rxbufstatus(1)) and (not spy_status_i.rxbufstatus(0)), -- 110
            count_o   => spy_mgt_buf_ovf
        );

    i_cnt_spy_mgt_buf_ovf_sync : xpm_cdc_gray
        generic map(
            DEST_SYNC_FF          => 4,
            REG_OUTPUT            => 0,
            WIDTH                 => 16
        )
        port map(
            src_clk      => spy_rx_usrclk_i,
            src_in_bin   => spy_mgt_buf_ovf,
            dest_clk     => clk_i,
            dest_out_bin => spy_mgt_buf_ovf_sync
        );
    
    -- elastic buffer underflow counter
    i_cnt_spy_mgt_buf_unf : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => spy_rx_usrclk_i,
            reset_i   => reset_i,
            en_i      => (spy_status_i.rxbufstatus(2)) and (not spy_status_i.rxbufstatus(1)) and (spy_status_i.rxbufstatus(0)), -- 101
            count_o   => spy_mgt_buf_unf
        );

    i_cnt_spy_mgt_buf_unf_sync : xpm_cdc_gray
        generic map(
            DEST_SYNC_FF          => 4,
            REG_OUTPUT            => 0,
            WIDTH                 => 16
        )
        port map(
            src_clk      => spy_rx_usrclk_i,
            src_in_bin   => spy_mgt_buf_unf,
            dest_clk     => clk_i,
            dest_out_bin => spy_mgt_buf_unf_sync
        );

    -- clock correction: idle word insertion counter 
    -- note: meaningful only for 1 GbE
    i_cnt_spy_clk_corr_add : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => spy_rx_usrclk_i,
            reset_i   => reset_i,
            en_i      => spy_status_i.rxclkcorcnt(1) and spy_status_i.rxclkcorcnt(0), -- 11
            count_o   => spy_clk_corr_add
        );

    i_cnt_spy_clk_corr_add_sync : xpm_cdc_gray
        generic map(
            DEST_SYNC_FF          => 4,
            REG_OUTPUT            => 0,
            WIDTH                 => 16
        )
        port map(
            src_clk      => spy_rx_usrclk_i,
            src_in_bin   => spy_clk_corr_add,
            dest_clk     => clk_i,
            dest_out_bin => spy_clk_corr_add_sync
        );

    -- clock correction: idle word drop counter 
    -- note: meaningful only for 1 GbE
    i_cnt_spy_clk_corr_drop : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => spy_rx_usrclk_i,
            reset_i   => reset_i,
            en_i      => spy_status_i.rxclkcorcnt(1) xor spy_status_i.rxclkcorcnt(0), -- 10 or 01
            count_o   => spy_clk_corr_drop
        );

    i_cnt_spy_clk_corr_drop_sync : xpm_cdc_gray
        generic map(
            DEST_SYNC_FF          => 4,
            REG_OUTPUT            => 0,
            WIDTH                 => 16
        )
        port map(
            src_clk      => spy_rx_usrclk_i,
            src_in_bin   => spy_clk_corr_drop,
            dest_clk     => clk_i,
            dest_out_bin => spy_clk_corr_drop_sync
        );

    -- not in table error counter
    -- note: meaningful only for 1 GbE
    i_cnt_spy_not_in_table : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => spy_rx_usrclk_i,
            reset_i   => reset_i,
            en_i      => spy_rx_data_i.rxnotintable(1) or spy_rx_data_i.rxnotintable(0),
            count_o   => spy_not_in_table
        );

    i_cnt_spy_not_in_table_sync : xpm_cdc_gray
        generic map(
            DEST_SYNC_FF          => 4,
            REG_OUTPUT            => 0,
            WIDTH                 => 16
        )
        port map(
            src_clk      => spy_rx_usrclk_i,
            src_in_bin   => spy_not_in_table,
            dest_clk     => clk_i,
            dest_out_bin => spy_not_in_table_sync
        );

    -- dispersion error counter
    -- note: meaningful only for 1 GbE
    i_cnt_spy_disperr : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => spy_rx_usrclk_i,
            reset_i   => reset_i,
            en_i      => spy_rx_data_i.rxdisperr(1) or spy_rx_data_i.rxdisperr(0),
            count_o   => spy_disperr
        );

    i_cnt_spy_disperr_sync : xpm_cdc_gray
        generic map(
            DEST_SYNC_FF          => 4,
            REG_OUTPUT            => 0,
            WIDTH                 => 16
        )
        port map(
            src_clk      => spy_rx_usrclk_i,
            src_in_bin   => spy_disperr,
            dest_clk     => clk_i,
            dest_out_bin => spy_disperr_sync
        );

    g_reg_ge11 : if g_GEM_STATION = 1 generate
    --==== Registers begin ge11 ==========================================================================
    --==== Registers end ge11 ============================================================================
    end generate;

    g_reg_ge21 : if g_GEM_STATION = 2 generate
    --==== Registers begin ge21 ==========================================================================
    --==== Registers end ge21 ============================================================================
    end generate;

    g_reg_me0 : if g_GEM_STATION = 0 generate
    --==== Registers begin me0 ==========================================================================
    --==== Registers end me0 ============================================================================
    end generate;
    
end oh_link_regs_arch;

