------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    12:22 2016-05-10
-- Module Name:    trigger
-- Description:    This module handles everything related to sbit cluster data (link synchronization, monitoring, local triggering, matching to L1A and reporting data to DAQ)  
------------------------------------------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

use work.common_pkg.all;
use work.csc_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity link_monitor is
    generic(
        g_NUM_OF_DMBs : integer
    );
    port(
        -- reset
        reset_i                 : in  std_logic;
        clk_i                   : in  std_logic;

        -- TTC
        ttc_clks_i              : in t_ttc_clks;
        ttc_cmds_i              : in t_ttc_cmds;

        -- DMB links
        csc_dmb_rx_usrclk_arr_i : in  std_logic_vector(g_NUM_OF_DMBs - 1 downto 0);
        csc_dmb_rx_data_arr_i   : in  t_mgt_16b_rx_data_arr(g_NUM_OF_DMBs - 1 downto 0);
        csc_dmb_rx_status_arr_i : in  t_mgt_status_arr(g_NUM_OF_DMBs - 1 downto 0);

        -- Spy link
        csc_spy_usrclk_i        : in  std_logic;
        csc_spy_rx_data_i       : in  t_mgt_16b_rx_data;
        csc_spy_rx_status_i     : in  t_mgt_status;
        
        -- IPbus
        ipb_reset_i             : in  std_logic;
        ipb_clk_i               : in  std_logic;
        ipb_miso_o              : out ipb_rbus;
        ipb_mosi_i              : in  ipb_wbus
    );
end link_monitor;

architecture link_monitor_arch of link_monitor is
    
    --=== resets ===--
    
    signal reset_global             : std_logic;
    signal reset_local              : std_logic;
    signal reset                    : std_logic;
    
    --=== counters ===--

    signal dmb_mgt_buf_ovf_arr      : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);
    signal dmb_mgt_buf_unf_arr      : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);
    signal dmb_not_in_table_arr     : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);
    signal dmb_disperr_arr          : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);
    signal dmb_clk_corr_add_arr     : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);
    signal dmb_clk_corr_drop_arr    : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);

    signal spy_mgt_buf_ovf          : std_logic_vector(15 downto 0);
    signal spy_mgt_buf_unf          : std_logic_vector(15 downto 0);
    signal spy_not_in_table         : std_logic_vector(15 downto 0);
    signal spy_disperr              : std_logic_vector(15 downto 0);
    signal spy_clk_corr_add         : std_logic_vector(15 downto 0);
    signal spy_clk_corr_drop        : std_logic_vector(15 downto 0);

    --=== Hard reset veto ===--
    constant HARD_RESET_VETO_TIME   : unsigned(23 downto 0) := x"b71b00"; -- number of 40MHz clock cycles to veto all counters after receiving a hard-reset TTC command
    signal hard_reset_countdown     : unsigned(23 downto 0) := HARD_RESET_VETO_TIME; -- countdown after receiving a hard reset 
    signal hard_reset_veto          : std_logic := '0';

    ------ Register signals begin (this section is generated by <csc_fed_repo_root>/scripts/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_LINKS_NUM_REGS - 1 downto 0);
    signal regs_write_arr       : t_std32_array(REG_LINKS_NUM_REGS - 1 downto 0);
    signal regs_addresses       : t_std32_array(REG_LINKS_NUM_REGS - 1 downto 0);
    signal regs_defaults        : t_std32_array(REG_LINKS_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_LINKS_NUM_REGS - 1 downto 0);
    signal regs_write_pulse_arr : std_logic_vector(REG_LINKS_NUM_REGS - 1 downto 0);
    signal regs_read_ready_arr  : std_logic_vector(REG_LINKS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_LINKS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_LINKS_NUM_REGS - 1 downto 0) := (others => '0');
    ------ Register signals end ----------------------------------------------
    
begin

    --================================--
    -- Resets  
    --================================--
    
    i_reset_sync : entity work.synch
        generic map(
            N_STAGES => 3
        )
        port map(
            async_i => reset_i,
            clk_i   => clk_i,
            sync_o  => reset_global
        );

    reset <= reset_global or reset_local;
    
    -- hard reset veto
    process(ttc_clks_i.clk_40)
    begin
        if (rising_edge(ttc_clks_i.clk_40)) then
            if (reset = '1') then
                hard_reset_countdown <= HARD_RESET_VETO_TIME;
                hard_reset_veto <= '1';
            else
                if (ttc_cmds_i.hard_reset = '1') then
                    hard_reset_countdown <= HARD_RESET_VETO_TIME;
                    hard_reset_veto <= '1';
                elsif (hard_reset_countdown = x"000000") then
                    hard_reset_countdown <= (others => '0');
                    hard_reset_veto <= '0';
                else
                    hard_reset_countdown <= hard_reset_countdown - 1;
                    hard_reset_veto <= '1';
                end if;
            end if;
        end if;
    end process;
    
    --================================--
    -- DMB link counetrs  
    --================================--
    
    i_dmbs : for i in 0 to g_NUM_OF_DMBs - 1 generate

        -- elastic buffer overflow counter
        i_cnt_dmb_mgt_buf_ovf : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => csc_dmb_rx_usrclk_arr_i(i),
                reset_i   => reset,
                en_i      => (csc_dmb_rx_status_arr_i(i).rxbufstatus(2)) and (csc_dmb_rx_status_arr_i(i).rxbufstatus(1)) and (not csc_dmb_rx_status_arr_i(i).rxbufstatus(0)) and not hard_reset_veto, -- 110
                count_o   => dmb_mgt_buf_ovf_arr(i)
            );
    
        -- elastic buffer underflow counter
        i_cnt_dmb_mgt_buf_unf : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => csc_dmb_rx_usrclk_arr_i(i),
                reset_i   => reset,
                en_i      => (csc_dmb_rx_status_arr_i(i).rxbufstatus(2)) and (not csc_dmb_rx_status_arr_i(i).rxbufstatus(1)) and (csc_dmb_rx_status_arr_i(i).rxbufstatus(0)) and not hard_reset_veto, -- 101
                count_o   => dmb_mgt_buf_unf_arr(i)
            );
    
        -- clock correction: idle word insertion counter 
        i_cnt_dmb_clk_corr_add : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => csc_dmb_rx_usrclk_arr_i(i),
                reset_i   => reset,
                en_i      => csc_dmb_rx_status_arr_i(i).rxclkcorcnt(1) and csc_dmb_rx_status_arr_i(i).rxclkcorcnt(0) and not hard_reset_veto, -- 11
                count_o   => dmb_clk_corr_add_arr(i)
            );
    
        -- clock correction: idle word drop counter 
        i_cnt_dmb_clk_corr_drop : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => csc_dmb_rx_usrclk_arr_i(i),
                reset_i   => reset,
                en_i      => (csc_dmb_rx_status_arr_i(i).rxclkcorcnt(1) xor csc_dmb_rx_status_arr_i(i).rxclkcorcnt(0)) and not hard_reset_veto, -- 10 or 01
                count_o   => dmb_clk_corr_drop_arr(i)
            );

        -- not in table error counter
        i_cnt_dmb_not_in_table : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => csc_dmb_rx_usrclk_arr_i(i),
                reset_i   => reset,
                en_i      => (csc_dmb_rx_data_arr_i(i).rxnotintable(1) or csc_dmb_rx_data_arr_i(i).rxnotintable(0)) and not hard_reset_veto,
                count_o   => dmb_not_in_table_arr(i)
            );

        -- disparity error counter
        i_cnt_dmb_disperr : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => csc_dmb_rx_usrclk_arr_i(i),
                reset_i   => reset,
                en_i      => (csc_dmb_rx_data_arr_i(i).rxdisperr(1) or csc_dmb_rx_data_arr_i(i).rxdisperr(0)) and not hard_reset_veto,
                count_o   => dmb_disperr_arr(i)
            );
      
    end generate i_dmbs;
    
    --================================--
    -- Spy link counters  
    --================================--

    -- elastic buffer overflow counter
    i_cnt_spy_mgt_buf_ovf : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => csc_spy_usrclk_i,
            reset_i   => reset,
            en_i      => (csc_spy_rx_status_i.rxbufstatus(2)) and (csc_spy_rx_status_i.rxbufstatus(1)) and (not csc_spy_rx_status_i.rxbufstatus(0)), -- 110
            count_o   => spy_mgt_buf_ovf
        );

    -- elastic buffer underflow counter
    i_cnt_spy_mgt_buf_unf : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => csc_spy_usrclk_i,
            reset_i   => reset,
            en_i      => (csc_spy_rx_status_i.rxbufstatus(2)) and (not csc_spy_rx_status_i.rxbufstatus(1)) and (csc_spy_rx_status_i.rxbufstatus(0)), -- 101
            count_o   => spy_mgt_buf_unf
        );

    -- clock correction: idle word insertion counter 
    i_cnt_spy_clk_corr_add : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => csc_spy_usrclk_i,
            reset_i   => reset,
            en_i      => csc_spy_rx_status_i.rxclkcorcnt(1) and csc_spy_rx_status_i.rxclkcorcnt(0), -- 11
            count_o   => spy_clk_corr_add
        );

    -- clock correction: idle word drop counter 
    i_cnt_spy_clk_corr_drop : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => csc_spy_usrclk_i,
            reset_i   => reset,
            en_i      => csc_spy_rx_status_i.rxclkcorcnt(1) xor csc_spy_rx_status_i.rxclkcorcnt(0), -- 10 or 01
            count_o   => spy_clk_corr_drop
        );

    -- not in table error counter
    i_cnt_spy_not_in_table : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => csc_spy_usrclk_i,
            reset_i   => reset,
            en_i      => csc_spy_rx_data_i.rxnotintable(1) or csc_spy_rx_data_i.rxnotintable(0),
            count_o   => spy_not_in_table
        );

    -- dispersion error counter
    i_cnt_dmb_disperr : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => csc_spy_usrclk_i,
            reset_i   => reset,
            en_i      => csc_spy_rx_data_i.rxdisperr(1) or csc_spy_rx_data_i.rxdisperr(0),
            count_o   => spy_disperr
        );
    
    --===============================================================================================
    -- this section is generated by <csc_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
           g_NUM_REGS             => REG_LINKS_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_LINKS_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_LINKS_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => ipb_clk_i,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => clk_i,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"000";
    regs_addresses(1)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"010";
    regs_addresses(2)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"011";
    regs_addresses(3)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"012";
    regs_addresses(4)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"020";
    regs_addresses(5)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"021";
    regs_addresses(6)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"022";
    regs_addresses(7)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"030";
    regs_addresses(8)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"031";
    regs_addresses(9)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"032";
    regs_addresses(10)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"040";
    regs_addresses(11)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"041";
    regs_addresses(12)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"042";
    regs_addresses(13)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"050";
    regs_addresses(14)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"051";
    regs_addresses(15)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"052";
    regs_addresses(16)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"060";
    regs_addresses(17)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"061";
    regs_addresses(18)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"062";
    regs_addresses(19)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"070";
    regs_addresses(20)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"071";
    regs_addresses(21)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"072";
    regs_addresses(22)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"080";
    regs_addresses(23)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"081";
    regs_addresses(24)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"082";
    regs_addresses(25)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"090";
    regs_addresses(26)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"091";
    regs_addresses(27)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"092";
    regs_addresses(28)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0a0";
    regs_addresses(29)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0a1";
    regs_addresses(30)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0a2";
    regs_addresses(31)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0b0";
    regs_addresses(32)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0b1";
    regs_addresses(33)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0b2";
    regs_addresses(34)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0c0";
    regs_addresses(35)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0c1";
    regs_addresses(36)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0c2";
    regs_addresses(37)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0d0";
    regs_addresses(38)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0d1";
    regs_addresses(39)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0d2";
    regs_addresses(40)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0e0";
    regs_addresses(41)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0e1";
    regs_addresses(42)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0e2";
    regs_addresses(43)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0f0";
    regs_addresses(44)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0f1";
    regs_addresses(45)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"0f2";
    regs_addresses(46)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"a00";
    regs_addresses(47)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"a01";
    regs_addresses(48)(REG_LINKS_ADDRESS_MSB downto REG_LINKS_ADDRESS_LSB) <= '0' & x"a02";

    -- Connect read signals
    regs_read_arr(1)(REG_LINKS_DMB0_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB0_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(0);
    regs_read_arr(1)(REG_LINKS_DMB0_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB0_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(0);
    regs_read_arr(2)(REG_LINKS_DMB0_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB0_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(0);
    regs_read_arr(2)(REG_LINKS_DMB0_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB0_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(0);
    regs_read_arr(3)(REG_LINKS_DMB0_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB0_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(0);
    regs_read_arr(3)(REG_LINKS_DMB0_DISPERR_CNT_MSB downto REG_LINKS_DMB0_DISPERR_CNT_LSB) <= dmb_disperr_arr(0);
    regs_read_arr(4)(REG_LINKS_DMB1_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB1_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(1);
    regs_read_arr(4)(REG_LINKS_DMB1_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB1_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(1);
    regs_read_arr(5)(REG_LINKS_DMB1_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB1_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(1);
    regs_read_arr(5)(REG_LINKS_DMB1_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB1_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(1);
    regs_read_arr(6)(REG_LINKS_DMB1_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB1_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(1);
    regs_read_arr(6)(REG_LINKS_DMB1_DISPERR_CNT_MSB downto REG_LINKS_DMB1_DISPERR_CNT_LSB) <= dmb_disperr_arr(1);
    regs_read_arr(7)(REG_LINKS_DMB2_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB2_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(2);
    regs_read_arr(7)(REG_LINKS_DMB2_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB2_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(2);
    regs_read_arr(8)(REG_LINKS_DMB2_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB2_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(2);
    regs_read_arr(8)(REG_LINKS_DMB2_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB2_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(2);
    regs_read_arr(9)(REG_LINKS_DMB2_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB2_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(2);
    regs_read_arr(9)(REG_LINKS_DMB2_DISPERR_CNT_MSB downto REG_LINKS_DMB2_DISPERR_CNT_LSB) <= dmb_disperr_arr(2);
    regs_read_arr(10)(REG_LINKS_DMB3_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB3_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(3);
    regs_read_arr(10)(REG_LINKS_DMB3_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB3_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(3);
    regs_read_arr(11)(REG_LINKS_DMB3_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB3_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(3);
    regs_read_arr(11)(REG_LINKS_DMB3_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB3_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(3);
    regs_read_arr(12)(REG_LINKS_DMB3_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB3_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(3);
    regs_read_arr(12)(REG_LINKS_DMB3_DISPERR_CNT_MSB downto REG_LINKS_DMB3_DISPERR_CNT_LSB) <= dmb_disperr_arr(3);
    regs_read_arr(13)(REG_LINKS_DMB4_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB4_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(4);
    regs_read_arr(13)(REG_LINKS_DMB4_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB4_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(4);
    regs_read_arr(14)(REG_LINKS_DMB4_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB4_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(4);
    regs_read_arr(14)(REG_LINKS_DMB4_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB4_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(4);
    regs_read_arr(15)(REG_LINKS_DMB4_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB4_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(4);
    regs_read_arr(15)(REG_LINKS_DMB4_DISPERR_CNT_MSB downto REG_LINKS_DMB4_DISPERR_CNT_LSB) <= dmb_disperr_arr(4);
    regs_read_arr(16)(REG_LINKS_DMB5_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB5_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(5);
    regs_read_arr(16)(REG_LINKS_DMB5_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB5_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(5);
    regs_read_arr(17)(REG_LINKS_DMB5_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB5_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(5);
    regs_read_arr(17)(REG_LINKS_DMB5_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB5_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(5);
    regs_read_arr(18)(REG_LINKS_DMB5_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB5_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(5);
    regs_read_arr(18)(REG_LINKS_DMB5_DISPERR_CNT_MSB downto REG_LINKS_DMB5_DISPERR_CNT_LSB) <= dmb_disperr_arr(5);
    regs_read_arr(19)(REG_LINKS_DMB6_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB6_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(6);
    regs_read_arr(19)(REG_LINKS_DMB6_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB6_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(6);
    regs_read_arr(20)(REG_LINKS_DMB6_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB6_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(6);
    regs_read_arr(20)(REG_LINKS_DMB6_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB6_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(6);
    regs_read_arr(21)(REG_LINKS_DMB6_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB6_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(6);
    regs_read_arr(21)(REG_LINKS_DMB6_DISPERR_CNT_MSB downto REG_LINKS_DMB6_DISPERR_CNT_LSB) <= dmb_disperr_arr(6);
    regs_read_arr(22)(REG_LINKS_DMB7_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB7_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(7);
    regs_read_arr(22)(REG_LINKS_DMB7_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB7_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(7);
    regs_read_arr(23)(REG_LINKS_DMB7_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB7_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(7);
    regs_read_arr(23)(REG_LINKS_DMB7_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB7_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(7);
    regs_read_arr(24)(REG_LINKS_DMB7_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB7_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(7);
    regs_read_arr(24)(REG_LINKS_DMB7_DISPERR_CNT_MSB downto REG_LINKS_DMB7_DISPERR_CNT_LSB) <= dmb_disperr_arr(7);
    regs_read_arr(25)(REG_LINKS_DMB8_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB8_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(8);
    regs_read_arr(25)(REG_LINKS_DMB8_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB8_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(8);
    regs_read_arr(26)(REG_LINKS_DMB8_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB8_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(8);
    regs_read_arr(26)(REG_LINKS_DMB8_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB8_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(8);
    regs_read_arr(27)(REG_LINKS_DMB8_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB8_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(8);
    regs_read_arr(27)(REG_LINKS_DMB8_DISPERR_CNT_MSB downto REG_LINKS_DMB8_DISPERR_CNT_LSB) <= dmb_disperr_arr(8);
    regs_read_arr(28)(REG_LINKS_DMB9_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB9_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(9);
    regs_read_arr(28)(REG_LINKS_DMB9_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB9_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(9);
    regs_read_arr(29)(REG_LINKS_DMB9_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB9_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(9);
    regs_read_arr(29)(REG_LINKS_DMB9_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB9_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(9);
    regs_read_arr(30)(REG_LINKS_DMB9_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB9_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(9);
    regs_read_arr(30)(REG_LINKS_DMB9_DISPERR_CNT_MSB downto REG_LINKS_DMB9_DISPERR_CNT_LSB) <= dmb_disperr_arr(9);
    regs_read_arr(31)(REG_LINKS_DMB10_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB10_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(10);
    regs_read_arr(31)(REG_LINKS_DMB10_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB10_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(10);
    regs_read_arr(32)(REG_LINKS_DMB10_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB10_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(10);
    regs_read_arr(32)(REG_LINKS_DMB10_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB10_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(10);
    regs_read_arr(33)(REG_LINKS_DMB10_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB10_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(10);
    regs_read_arr(33)(REG_LINKS_DMB10_DISPERR_CNT_MSB downto REG_LINKS_DMB10_DISPERR_CNT_LSB) <= dmb_disperr_arr(10);
    regs_read_arr(34)(REG_LINKS_DMB11_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB11_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(11);
    regs_read_arr(34)(REG_LINKS_DMB11_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB11_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(11);
    regs_read_arr(35)(REG_LINKS_DMB11_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB11_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(11);
    regs_read_arr(35)(REG_LINKS_DMB11_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB11_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(11);
    regs_read_arr(36)(REG_LINKS_DMB11_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB11_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(11);
    regs_read_arr(36)(REG_LINKS_DMB11_DISPERR_CNT_MSB downto REG_LINKS_DMB11_DISPERR_CNT_LSB) <= dmb_disperr_arr(11);
    regs_read_arr(37)(REG_LINKS_DMB12_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB12_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(12);
    regs_read_arr(37)(REG_LINKS_DMB12_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB12_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(12);
    regs_read_arr(38)(REG_LINKS_DMB12_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB12_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(12);
    regs_read_arr(38)(REG_LINKS_DMB12_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB12_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(12);
    regs_read_arr(39)(REG_LINKS_DMB12_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB12_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(12);
    regs_read_arr(39)(REG_LINKS_DMB12_DISPERR_CNT_MSB downto REG_LINKS_DMB12_DISPERR_CNT_LSB) <= dmb_disperr_arr(12);
    regs_read_arr(40)(REG_LINKS_DMB13_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB13_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(13);
    regs_read_arr(40)(REG_LINKS_DMB13_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB13_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(13);
    regs_read_arr(41)(REG_LINKS_DMB13_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB13_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(13);
    regs_read_arr(41)(REG_LINKS_DMB13_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB13_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(13);
    regs_read_arr(42)(REG_LINKS_DMB13_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB13_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(13);
    regs_read_arr(42)(REG_LINKS_DMB13_DISPERR_CNT_MSB downto REG_LINKS_DMB13_DISPERR_CNT_LSB) <= dmb_disperr_arr(13);
    regs_read_arr(43)(REG_LINKS_DMB14_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_DMB14_MGT_BUF_OVF_CNT_LSB) <= dmb_mgt_buf_ovf_arr(14);
    regs_read_arr(43)(REG_LINKS_DMB14_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_DMB14_MGT_BUF_UNF_CNT_LSB) <= dmb_mgt_buf_unf_arr(14);
    regs_read_arr(44)(REG_LINKS_DMB14_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_DMB14_CLK_CORR_ADD_CNT_LSB) <= dmb_clk_corr_add_arr(14);
    regs_read_arr(44)(REG_LINKS_DMB14_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_DMB14_CLK_CORR_DROP_CNT_LSB) <= dmb_clk_corr_drop_arr(14);
    regs_read_arr(45)(REG_LINKS_DMB14_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_DMB14_NOT_IN_TABLE_CNT_LSB) <= dmb_not_in_table_arr(14);
    regs_read_arr(45)(REG_LINKS_DMB14_DISPERR_CNT_MSB downto REG_LINKS_DMB14_DISPERR_CNT_LSB) <= dmb_disperr_arr(14);
    regs_read_arr(46)(REG_LINKS_SPY_MGT_BUF_OVF_CNT_MSB downto REG_LINKS_SPY_MGT_BUF_OVF_CNT_LSB) <= spy_mgt_buf_ovf;
    regs_read_arr(46)(REG_LINKS_SPY_MGT_BUF_UNF_CNT_MSB downto REG_LINKS_SPY_MGT_BUF_UNF_CNT_LSB) <= spy_mgt_buf_unf;
    regs_read_arr(47)(REG_LINKS_SPY_CLK_CORR_ADD_CNT_MSB downto REG_LINKS_SPY_CLK_CORR_ADD_CNT_LSB) <= spy_clk_corr_add;
    regs_read_arr(47)(REG_LINKS_SPY_CLK_CORR_DROP_CNT_MSB downto REG_LINKS_SPY_CLK_CORR_DROP_CNT_LSB) <= spy_clk_corr_drop;
    regs_read_arr(48)(REG_LINKS_SPY_NOT_IN_TABLE_CNT_MSB downto REG_LINKS_SPY_NOT_IN_TABLE_CNT_LSB) <= spy_not_in_table;
    regs_read_arr(48)(REG_LINKS_SPY_DISPERR_CNT_MSB downto REG_LINKS_SPY_DISPERR_CNT_LSB) <= spy_disperr;

    -- Connect write signals

    -- Connect write pulse signals
    reset_local <= regs_write_pulse_arr(0);

    -- Connect write done signals

    -- Connect read pulse signals

    -- Connect read ready signals

    -- Defaults

    -- Define writable regs

    --==== Registers end ============================================================================
    
end link_monitor_arch;

