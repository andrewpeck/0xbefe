library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package project_config is
    

end package project_config;

