------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    12:22 2016-05-10
-- Module Name:    trigger
-- Description:    This module handles everything related to sbit cluster data (link synchronization, monitoring, local triggering, matching to L1A and reporting data to DAQ)  
------------------------------------------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

use work.common_pkg.all;
use work.csc_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity link_monitor is
    generic(
        g_NUM_OF_DMBs       : integer;
        g_NUM_GBT_LINKS     : integer;
        g_IPB_CLK_PERIOD_NS : integer
    );
    port(
        -- reset
        reset_i                 : in  std_logic;
        clk_i                   : in  std_logic;

        -- TTC
        ttc_clks_i              : in t_ttc_clks;
        ttc_cmds_i              : in t_ttc_cmds;

        -- DMB links
        dmb_rx_usrclk_i         : in  std_logic;
        dmb_rx_data_arr_i       : in  t_mgt_16b_rx_data_arr(g_NUM_OF_DMBs - 1 downto 0);
        dmb_rx_status_arr_i     : in  t_mgt_status_arr(g_NUM_OF_DMBs - 1 downto 0);

        -- GBT links
        gbt_link_status_arr_i   : in t_gbt_link_status_arr(g_NUM_GBT_LINKS - 1 downto 0);

        -- Spy link
        spy_usrclk_i            : in  std_logic;
        spy_rx_data_i           : in  t_mgt_16b_rx_data;
        spy_rx_status_i         : in  t_mgt_status;
        
        -- IPbus
        ipb_reset_i             : in  std_logic;
        ipb_clk_i               : in  std_logic;
        ipb_miso_o              : out ipb_rbus;
        ipb_mosi_i              : in  ipb_wbus
    );
end link_monitor;

architecture link_monitor_arch of link_monitor is
    
    --=== resets ===--
    
    signal reset_global             : std_logic;
    signal reset_local              : std_logic;
    signal reset                    : std_logic;
    
    --=== counters ===--

    signal dmb_mgt_buf_ovf_arr      : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);
    signal dmb_mgt_buf_unf_arr      : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);
    signal dmb_not_in_table_arr     : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);
    signal dmb_disperr_arr          : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);
    signal dmb_clk_corr_add_arr     : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);
    signal dmb_clk_corr_drop_arr    : t_std16_array(g_NUM_OF_DMBs - 1 downto 0);

    signal spy_mgt_buf_ovf          : std_logic_vector(15 downto 0);
    signal spy_mgt_buf_unf          : std_logic_vector(15 downto 0);
    signal spy_not_in_table         : std_logic_vector(15 downto 0);
    signal spy_disperr              : std_logic_vector(15 downto 0);
    signal spy_clk_corr_add         : std_logic_vector(15 downto 0);
    signal spy_clk_corr_drop        : std_logic_vector(15 downto 0);

    --=== Hard reset veto ===--
    constant HARD_RESET_VETO_TIME   : unsigned(23 downto 0) := x"b71b00"; -- number of 40MHz clock cycles to veto all counters after receiving a hard-reset TTC command
    signal hard_reset_countdown     : unsigned(23 downto 0) := HARD_RESET_VETO_TIME; -- countdown after receiving a hard reset 
    signal hard_reset_veto          : std_logic := '0';

    ------ Register signals begin (this section is generated by <csc_fed_repo_root>/scripts/generate_registers.py -- do not edit)
    ------ Register signals end ----------------------------------------------
    
begin

    --================================--
    -- Resets  
    --================================--
    
    i_reset_sync : entity work.synch
        generic map(
            N_STAGES => 3
        )
        port map(
            async_i => reset_i,
            clk_i   => clk_i,
            sync_o  => reset_global
        );

    reset <= reset_global or reset_local;
    
    -- hard reset veto
    process(ttc_clks_i.clk_40)
    begin
        if (rising_edge(ttc_clks_i.clk_40)) then
            if (reset = '1') then
                hard_reset_countdown <= HARD_RESET_VETO_TIME;
                hard_reset_veto <= '1';
            else
                if (ttc_cmds_i.hard_reset = '1') then
                    hard_reset_countdown <= HARD_RESET_VETO_TIME;
                    hard_reset_veto <= '1';
                elsif (hard_reset_countdown = x"000000") then
                    hard_reset_countdown <= (others => '0');
                    hard_reset_veto <= '0';
                else
                    hard_reset_countdown <= hard_reset_countdown - 1;
                    hard_reset_veto <= '1';
                end if;
            end if;
        end if;
    end process;
    
    --================================--
    -- DMB link counetrs  
    --================================--
    
    i_dmbs : for i in 0 to g_NUM_OF_DMBs - 1 generate

        -- elastic buffer overflow counter
        i_cnt_dmb_mgt_buf_ovf : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => dmb_rx_usrclk_i,
                reset_i   => reset,
                en_i      => (dmb_rx_status_arr_i(i).rxbufstatus(2)) and (dmb_rx_status_arr_i(i).rxbufstatus(1)) and (not dmb_rx_status_arr_i(i).rxbufstatus(0)) and not hard_reset_veto, -- 110
                count_o   => dmb_mgt_buf_ovf_arr(i)
            );
    
        -- elastic buffer underflow counter
        i_cnt_dmb_mgt_buf_unf : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => dmb_rx_usrclk_i,
                reset_i   => reset,
                en_i      => (dmb_rx_status_arr_i(i).rxbufstatus(2)) and (not dmb_rx_status_arr_i(i).rxbufstatus(1)) and (dmb_rx_status_arr_i(i).rxbufstatus(0)) and not hard_reset_veto, -- 101
                count_o   => dmb_mgt_buf_unf_arr(i)
            );
    
        -- clock correction: idle word insertion counter 
        i_cnt_dmb_clk_corr_add : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => dmb_rx_usrclk_i,
                reset_i   => reset,
                en_i      => dmb_rx_status_arr_i(i).rxclkcorcnt(1) and dmb_rx_status_arr_i(i).rxclkcorcnt(0) and not hard_reset_veto, -- 11
                count_o   => dmb_clk_corr_add_arr(i)
            );
    
        -- clock correction: idle word drop counter 
        i_cnt_dmb_clk_corr_drop : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => dmb_rx_usrclk_i,
                reset_i   => reset,
                en_i      => (dmb_rx_status_arr_i(i).rxclkcorcnt(1) xor dmb_rx_status_arr_i(i).rxclkcorcnt(0)) and not hard_reset_veto, -- 10 or 01
                count_o   => dmb_clk_corr_drop_arr(i)
            );

        -- not in table error counter
        i_cnt_dmb_not_in_table : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => dmb_rx_usrclk_i,
                reset_i   => reset,
                en_i      => (dmb_rx_data_arr_i(i).rxnotintable(1) or dmb_rx_data_arr_i(i).rxnotintable(0)) and not hard_reset_veto,
                count_o   => dmb_not_in_table_arr(i)
            );

        -- disparity error counter
        i_cnt_dmb_disperr : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 16
            )
            port map(
                ref_clk_i => dmb_rx_usrclk_i,
                reset_i   => reset,
                en_i      => (dmb_rx_data_arr_i(i).rxdisperr(1) or dmb_rx_data_arr_i(i).rxdisperr(0)) and not hard_reset_veto,
                count_o   => dmb_disperr_arr(i)
            );
      
    end generate i_dmbs;
    
    --================================--
    -- Spy link counters  
    --================================--

    -- elastic buffer overflow counter
    i_cnt_spy_mgt_buf_ovf : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => spy_usrclk_i,
            reset_i   => reset,
            en_i      => (spy_rx_status_i.rxbufstatus(2)) and (spy_rx_status_i.rxbufstatus(1)) and (not spy_rx_status_i.rxbufstatus(0)), -- 110
            count_o   => spy_mgt_buf_ovf
        );

    -- elastic buffer underflow counter
    i_cnt_spy_mgt_buf_unf : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => spy_usrclk_i,
            reset_i   => reset,
            en_i      => (spy_rx_status_i.rxbufstatus(2)) and (not spy_rx_status_i.rxbufstatus(1)) and (spy_rx_status_i.rxbufstatus(0)), -- 101
            count_o   => spy_mgt_buf_unf
        );

    -- clock correction: idle word insertion counter 
    i_cnt_spy_clk_corr_add : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => spy_usrclk_i,
            reset_i   => reset,
            en_i      => spy_rx_status_i.rxclkcorcnt(1) and spy_rx_status_i.rxclkcorcnt(0), -- 11
            count_o   => spy_clk_corr_add
        );

    -- clock correction: idle word drop counter 
    i_cnt_spy_clk_corr_drop : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => spy_usrclk_i,
            reset_i   => reset,
            en_i      => spy_rx_status_i.rxclkcorcnt(1) xor spy_rx_status_i.rxclkcorcnt(0), -- 10 or 01
            count_o   => spy_clk_corr_drop
        );

    -- not in table error counter
    i_cnt_spy_not_in_table : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => spy_usrclk_i,
            reset_i   => reset,
            en_i      => spy_rx_data_i.rxnotintable(1) or spy_rx_data_i.rxnotintable(0),
            count_o   => spy_not_in_table
        );

    -- dispersion error counter
    i_cnt_dmb_disperr : entity work.counter
        generic map(
            g_COUNTER_WIDTH => 16
        )
        port map(
            ref_clk_i => spy_usrclk_i,
            reset_i   => reset,
            en_i      => spy_rx_data_i.rxdisperr(1) or spy_rx_data_i.rxdisperr(0),
            count_o   => spy_disperr
        );
    
    --===============================================================================================
    -- this section is generated by <csc_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    --==== Registers end ============================================================================
    
end link_monitor_arch;

