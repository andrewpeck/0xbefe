------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    2020-07-16
-- Module Name:    GEM_LOADER
-- Description:    This module implements the so called gemloader module which stores the frontend firmware, and streams it to the gem logic on request.
--                 This version uses a QDR II+ chip for storing the bitfile (this was written for CTP7 that has CY7C1263KV18)
------------------------------------------------------------------------------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library UNISIM;
use UNISIM.VComponents.all;

use work.ttc_pkg.all;
use work.common_pkg.all;
use work.gem_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity promless is
    port (
        reset_i             : in  std_logic;
        
        -- QDR interface
        qdriip_cq_p_i       : in  std_logic;
        qdriip_cq_n_i       : in  std_logic;
        qdriip_q_i          : in  std_logic_vector(17 downto 0);
        qdriip_k_p_o        : out std_logic;
        qdriip_k_n_o        : out std_logic;
        qdriip_d_o          : out std_logic_vector(17 downto 0);
        qdriip_sa_o         : out std_logic_vector(18 downto 0);
        qdriip_w_n_o        : out std_logic;
        qdriip_r_n_o        : out std_logic;
        qdriip_bw_n_o       : out std_logic_vector(1 downto 0);
        qdriip_dll_off_n_o  : out std_logic;        
        
        -- user interface
        clk40_i             : in  std_logic;
        to_gem_loader_i     : in  t_to_gem_loader;
        from_gem_loader_o   : out t_from_gem_loader;        
        
        -- IPbus
        ipb_reset_i         : in  std_logic;
        ipb_clk_i           : in  std_logic;
        ipb_miso_o          : out ipb_rbus;
        ipb_mosi_i          : in  ipb_wbus                
    );
end promless;

architecture promless_arch of promless is

    signal qdr_k_clk        : std_logic;
    signal qdr_cq_clk       : std_logic;
    signal qdr_q            : std_logic_vector(35 downto 0);
    signal qdr_d            : std_logic_vector(35 downto 0);

    type t_qdr_state is (IDLE, WRITE1, WRITE2, READ_WAIT, READ1, READ2);

    signal qdr_write_data   : std_logic_vector(17 downto 0);
    signal qdr_read_data    : std_logic_vector(71 downto 0);
    
    -- slow control signals
    signal sc_write_addr    : std_logic_vector(18 downto 0);
    signal sc_read_addr     : std_logic_vector(18 downto 0);
    signal sc_qdr_addr      : std_logic_vector(18 downto 0);
    signal sc_write_req     : std_logic;
    signal sc_read_req      : std_logic;
    signal sc_addr_reset    : std_logic;
    signal sc_bw            : std_logic_vector(3 downto 0);
    signal sc_wps           : std_logic;
    signal sc_rps           : std_logic;
    
    -- streaming signals
    signal streaming_mode   : std_logic;
    
    signal st_rps           : std_logic;
    signal st_addr          : std_logic_vector(18 downto 0);

    ------ Register signals begin (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    ------ Register signals end ----------------------------------------------
        
begin

    -- I/O buffers

    qdr_k_clk <= clk40_i;
    qdriip_dll_off_n_o <= '0'; -- turn off the PLL on the chip, and use it in QDR I mode
    qdriip_sa_o <= sc_qdr_addr when streaming_mode = '0' else st_addr;
    qdriip_w_n_o <= not sc_wps when streaming_mode = '0' else '1';
    qdriip_r_n_o <= not sc_rps when streaming_mode = '0' else st_rps;

    i_cq_clk_ibuf : IBUFGDS
        generic map(
            DIFF_TERM        => true,
            IBUF_LOW_PWR     => false
        )
        port map(
            O  => qdr_cq_clk,
            I  => qdriip_cq_p_i,
            IB => qdriip_cq_n_i
        );

    i_k_clk_obuf : OBUFDS
        port map(
            O  => qdriip_k_p_o,
            OB => qdriip_k_n_o,
            I  => qdr_k_clk
        );

    g_data_bus_buf: for i in 0 to 17 generate
        i_q_iddr : IDDR
            generic map(
                DDR_CLK_EDGE => "SAME_EDGE"
            )
            port map(
                q1 => qdr_q(i),
                q2 => qdr_q(i+18),
                c  => qdr_cq_clk,
                ce => '1',
                d  => qdriip_q_i(i),
                r  => '0',
                s  => '0'
            );    
    
        i_d_oddr : ODDR
            generic map(
                DDR_CLK_EDGE => "SAME_EDGE"
            )
            port map(
                q  => qdriip_d_o(i),
                c  => qdr_k_clk,
                ce => '1',
                d1 => qdr_d(i),
                d2 => qdr_d(i+18),
                r  => '0',
                s  => '0'
            );
    end generate;

    g_bw_buf: for i in 0 to 1 generate
        i_bw_oddr : ODDR
            generic map(
                DDR_CLK_EDGE => "SAME_EDGE"
            )
            port map(
                q  => qdriip_bw_n_o(i),
                c  => qdr_k_clk,
                ce => '1',
                d1 => not qdr_bw(i),
                d2 => not qdr_bw(i+2),
                r  => '0',
                s  => '0'
            );
    end generate;

    process (qdr_k_clk)
    begin
        if rising_edge(qdr_k_clk) then
            if (reset_i = '1' or sc_addr_reset = '1') then
                sc_write_addr <= (others => '0');
                sc_read_addr <= (others => '0');
                sc_qdr_addr <= (others => '0');
                sc_bw <= (others => '0');
                sc_wps <= '0';
                sc_rps <= '0';
            else
                if (sc_write_req = '1') then
                    sc_qdr_addr <= sc_write_addr;
                    -- ok, dropped it at this point since we seem to have gotten gemloader to work.. can pick it up here at a later date
                else
                end if;
            end if;
        end if;
    end process;

    --===============================================================================================
    -- this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    --==== Registers end ============================================================================
    
end promless_arch;
