------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    2020-06-16
-- Module Name:    MGT_SLOW_CONTROL 
-- Description:    Slow control interface for MGTs    
------------------------------------------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_misc.all;

library unisim;
use unisim.vcomponents.all;

library xpm;
use xpm.vcomponents.all;

use work.common_pkg.all;
use work.mgt_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity mgt_slow_control is
    generic(
        g_NUM_CHANNELS          : integer
    );
    port(
        
        clk_stable_i            : in  std_logic;
        
        mgt_clks_arr_i          : in  t_mgt_clk_in_arr(g_NUM_CHANNELS - 1 downto 0);

        tx_reset_arr_o          : out std_logic_vector(g_NUM_CHANNELS - 1 downto 0);
        rx_reset_arr_o          : out std_logic_vector(g_NUM_CHANNELS - 1 downto 0);
        
        tx_slow_ctrl_arr_o      : out t_mgt_tx_slow_ctrl_arr(g_NUM_CHANNELS - 1 downto 0);
        rx_slow_ctrl_arr_o      : out t_mgt_rx_slow_ctrl_arr(g_NUM_CHANNELS - 1 downto 0);
        misc_ctrl_arr_o         : out t_mgt_misc_ctrl_arr(g_NUM_CHANNELS - 1 downto 0);

        tx_status_arr_i         : in  t_mgt_tx_status_arr(g_NUM_CHANNELS - 1 downto 0);
        rx_status_arr_i         : in  t_mgt_rx_status_arr(g_NUM_CHANNELS - 1 downto 0);
        misc_status_arr_i       : in  t_mgt_misc_status_arr(g_NUM_CHANNELS - 1 downto 0);
        ibert_eyescanreset_i    : in  std_logic_vector(g_NUM_CHANNELS - 1 downto 0);
        
        tx_reset_done_arr_i     : in  std_logic_vector(g_NUM_CHANNELS - 1 downto 0);
        rx_reset_done_arr_i     : in  std_logic_vector(g_NUM_CHANNELS - 1 downto 0);
        tx_phalign_done_arr_i   : in  std_logic_vector(g_NUM_CHANNELS - 1 downto 0);
        rx_phalign_done_arr_i   : in  std_logic_vector(g_NUM_CHANNELS - 1 downto 0);
        
        cpll_status_arr_i       : in  t_mgt_cpll_status_arr(g_NUM_CHANNELS - 1 downto 0);
        
        ipb_clk_i               : in  std_logic;
        ipb_reset_i             : in  std_logic;
        ipb_mosi_i              : in  ipb_wbus;
        ipb_miso_o              : out ipb_rbus
    );
end mgt_slow_control;

architecture mgt_slow_control_arch of mgt_slow_control is

    signal tx_slow_ctrl_arr         : t_mgt_tx_slow_ctrl_arr(g_NUM_CHANNELS - 1 downto 0);
    signal rx_slow_ctrl_arr         : t_mgt_rx_slow_ctrl_arr(g_NUM_CHANNELS - 1 downto 0);
    signal misc_ctrl_arr            : t_mgt_misc_ctrl_arr(g_NUM_CHANNELS - 1 downto 0);

    signal reset_arr                : std_logic_vector(g_NUM_CHANNELS - 1 downto 0);
    signal loopback_arr             : std_logic_vector(g_NUM_CHANNELS - 1 downto 0);
    signal txpd_arr                 : std_logic_vector(g_NUM_CHANNELS - 1 downto 0);
    signal rxpd_arr                 : std_logic_vector(g_NUM_CHANNELS - 1 downto 0);
    signal prbs_err_reset_arr       : std_logic_vector(g_NUM_CHANNELS - 1 downto 0);
    signal prbs_err_reset_sync_arr  : std_logic_vector(g_NUM_CHANNELS - 1 downto 0);    
    signal prbs_err_cnt_arr         : t_std32_array(g_NUM_CHANNELS - 1 downto 0);    
    signal prbs_err_cnt_sync_arr    : t_std32_array(g_NUM_CHANNELS - 1 downto 0);    

    ------ Register signals begin (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_OPTICAL_LINKS_NUM_REGS - 1 downto 0);
    signal regs_write_arr       : t_std32_array(REG_OPTICAL_LINKS_NUM_REGS - 1 downto 0);
    signal regs_addresses       : t_std32_array(REG_OPTICAL_LINKS_NUM_REGS - 1 downto 0);
    signal regs_defaults        : t_std32_array(REG_OPTICAL_LINKS_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_OPTICAL_LINKS_NUM_REGS - 1 downto 0);
    signal regs_write_pulse_arr : std_logic_vector(REG_OPTICAL_LINKS_NUM_REGS - 1 downto 0);
    signal regs_read_ready_arr  : std_logic_vector(REG_OPTICAL_LINKS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_OPTICAL_LINKS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_OPTICAL_LINKS_NUM_REGS - 1 downto 0) := (others => '0');
    ------ Register signals end ----------------------------------------------

begin

    tx_reset_arr_o <= reset_arr;
    rx_reset_arr_o <= reset_arr;
    
    tx_slow_ctrl_arr_o <= tx_slow_ctrl_arr;
    rx_slow_ctrl_arr_o <= rx_slow_ctrl_arr;
    misc_ctrl_arr_o <= misc_ctrl_arr;
    
    g_channels : for chan in 0 to g_NUM_CHANNELS - 1 generate
        -- ibert
        misc_ctrl_arr(chan).eyescanreset <= ibert_eyescanreset_i(chan);
    
        -- loopback and PD controll
        misc_ctrl_arr(chan).loopback <= "000" when loopback_arr(chan) = '0' else "010";
        tx_slow_ctrl_arr(chan).txpd <= "00" when txpd_arr(chan) = '0' else "11";
        rx_slow_ctrl_arr(chan).rxpd <= "00" when rxpd_arr(chan) = '0' else "11";
        rx_slow_ctrl_arr(chan).rxbufreset <= '0';

        -- prbs error counting
        i_sync_prbs_err_reset : entity work.synch generic map(N_STAGES => 3, IS_RESET => false) port map(async_i => prbs_err_reset_arr(chan), clk_i => mgt_clks_arr_i(chan).rxusrclk2, sync_o  => prbs_err_reset_sync_arr(chan));        
        i_prbs_cnt : entity work.counter
            generic map(
                g_COUNTER_WIDTH  => 32,
                g_ALLOW_ROLLOVER => false
            )
            port map(
                ref_clk_i => mgt_clks_arr_i(chan).rxusrclk2,
                reset_i   => prbs_err_reset_sync_arr(chan),
                en_i      => rx_status_arr_i(chan).rxprbserr,
                count_o   => prbs_err_cnt_arr(chan)
            );
        
        i_sync_prbs_err_cnt : xpm_cdc_gray
            generic map(
                DEST_SYNC_FF          => 2,
                WIDTH                 => 32
            )
            port map(
                src_clk      => mgt_clks_arr_i(chan).rxusrclk2,
                src_in_bin   => prbs_err_cnt_arr(chan),
                dest_clk     => clk_stable_i,
                dest_out_bin => prbs_err_cnt_sync_arr(chan)
            );
        
    end generate;

    --===============================================================================================
    -- this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
           g_NUM_REGS             => REG_OPTICAL_LINKS_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_OPTICAL_LINKS_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_OPTICAL_LINKS_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => ipb_clk_i,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => clk_stable_i,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0000";
    regs_addresses(1)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0001";
    regs_addresses(2)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0002";
    regs_addresses(3)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0003";
    regs_addresses(4)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0004";
    regs_addresses(5)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0005";
    regs_addresses(6)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0020";
    regs_addresses(7)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0021";
    regs_addresses(8)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0040";
    regs_addresses(9)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0041";
    regs_addresses(10)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0042";
    regs_addresses(11)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0043";
    regs_addresses(12)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0044";
    regs_addresses(13)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0045";
    regs_addresses(14)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0060";
    regs_addresses(15)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0061";
    regs_addresses(16)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0080";
    regs_addresses(17)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0081";
    regs_addresses(18)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0082";
    regs_addresses(19)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0083";
    regs_addresses(20)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0084";
    regs_addresses(21)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0085";
    regs_addresses(22)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"00a0";
    regs_addresses(23)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"00a1";
    regs_addresses(24)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"00c0";
    regs_addresses(25)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"00c1";
    regs_addresses(26)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"00c2";
    regs_addresses(27)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"00c3";
    regs_addresses(28)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"00c4";
    regs_addresses(29)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"00c5";
    regs_addresses(30)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"00e0";
    regs_addresses(31)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"00e1";
    regs_addresses(32)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0100";
    regs_addresses(33)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0101";
    regs_addresses(34)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0102";
    regs_addresses(35)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0103";
    regs_addresses(36)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0104";
    regs_addresses(37)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0105";
    regs_addresses(38)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0120";
    regs_addresses(39)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0121";
    regs_addresses(40)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0140";
    regs_addresses(41)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0141";
    regs_addresses(42)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0142";
    regs_addresses(43)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0143";
    regs_addresses(44)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0144";
    regs_addresses(45)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0145";
    regs_addresses(46)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0160";
    regs_addresses(47)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0161";
    regs_addresses(48)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0180";
    regs_addresses(49)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0181";
    regs_addresses(50)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0182";
    regs_addresses(51)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0183";
    regs_addresses(52)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0184";
    regs_addresses(53)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0185";
    regs_addresses(54)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"01a0";
    regs_addresses(55)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"01a1";
    regs_addresses(56)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"01c0";
    regs_addresses(57)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"01c1";
    regs_addresses(58)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"01c2";
    regs_addresses(59)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"01c3";
    regs_addresses(60)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"01c4";
    regs_addresses(61)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"01c5";
    regs_addresses(62)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"01e0";
    regs_addresses(63)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"01e1";
    regs_addresses(64)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0200";
    regs_addresses(65)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0201";
    regs_addresses(66)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0202";
    regs_addresses(67)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0203";
    regs_addresses(68)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0204";
    regs_addresses(69)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0205";
    regs_addresses(70)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0220";
    regs_addresses(71)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0221";
    regs_addresses(72)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0240";
    regs_addresses(73)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0241";
    regs_addresses(74)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0242";
    regs_addresses(75)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0243";
    regs_addresses(76)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0244";
    regs_addresses(77)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0245";
    regs_addresses(78)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0260";
    regs_addresses(79)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0261";
    regs_addresses(80)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0280";
    regs_addresses(81)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0281";
    regs_addresses(82)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0282";
    regs_addresses(83)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0283";
    regs_addresses(84)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0284";
    regs_addresses(85)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0285";
    regs_addresses(86)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"02a0";
    regs_addresses(87)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"02a1";
    regs_addresses(88)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"02c0";
    regs_addresses(89)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"02c1";
    regs_addresses(90)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"02c2";
    regs_addresses(91)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"02c3";
    regs_addresses(92)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"02c4";
    regs_addresses(93)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"02c5";
    regs_addresses(94)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"02e0";
    regs_addresses(95)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"02e1";
    regs_addresses(96)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0300";
    regs_addresses(97)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0301";
    regs_addresses(98)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0302";
    regs_addresses(99)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0303";
    regs_addresses(100)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0304";
    regs_addresses(101)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0305";
    regs_addresses(102)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0320";
    regs_addresses(103)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0321";
    regs_addresses(104)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0340";
    regs_addresses(105)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0341";
    regs_addresses(106)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0342";
    regs_addresses(107)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0343";
    regs_addresses(108)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0344";
    regs_addresses(109)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0345";
    regs_addresses(110)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0360";
    regs_addresses(111)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0361";
    regs_addresses(112)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0380";
    regs_addresses(113)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0381";
    regs_addresses(114)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0382";
    regs_addresses(115)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0383";
    regs_addresses(116)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0384";
    regs_addresses(117)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"0385";
    regs_addresses(118)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"03a0";
    regs_addresses(119)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"03a1";
    regs_addresses(120)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"03c0";
    regs_addresses(121)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"03c1";
    regs_addresses(122)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"03c2";
    regs_addresses(123)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"03c3";
    regs_addresses(124)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"03c4";
    regs_addresses(125)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"03c5";
    regs_addresses(126)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"03e0";
    regs_addresses(127)(REG_OPTICAL_LINKS_ADDRESS_MSB downto REG_OPTICAL_LINKS_ADDRESS_LSB) <= x"03e1";

    -- Connect read signals
    regs_read_arr(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(0);
    regs_read_arr(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(0);
    regs_read_arr(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(0).txpolarity;
    regs_read_arr(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(0).rxpolarity;
    regs_read_arr(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_LOOPBACK_BIT) <= loopback_arr(0);
    regs_read_arr(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(0).txinhibit;
    regs_read_arr(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(0).rxlpmen;
    regs_read_arr(2)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(0).txdiffctrl;
    regs_read_arr(2)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(0).txprecursor;
    regs_read_arr(2)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(0).txpostcursor;
    regs_read_arr(2)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(0).txmaincursor;
    regs_read_arr(3)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(0).rxprbssel;
    regs_read_arr(3)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(0).txprbssel;
    regs_read_arr(6)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(0);
    regs_read_arr(6)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(0);
    regs_read_arr(6)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(0);
    regs_read_arr(6)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(0);
    regs_read_arr(6)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(0).powergood;
    regs_read_arr(6)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(0).cplllock;
    regs_read_arr(6)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(0).cpllrefclklost;
    regs_read_arr(7)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(0);
    regs_read_arr(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(1);
    regs_read_arr(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(1);
    regs_read_arr(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(1).txpolarity;
    regs_read_arr(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(1).rxpolarity;
    regs_read_arr(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_LOOPBACK_BIT) <= loopback_arr(1);
    regs_read_arr(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(1).txinhibit;
    regs_read_arr(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(1).rxlpmen;
    regs_read_arr(10)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(1).txdiffctrl;
    regs_read_arr(10)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(1).txprecursor;
    regs_read_arr(10)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(1).txpostcursor;
    regs_read_arr(10)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(1).txmaincursor;
    regs_read_arr(11)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(1).rxprbssel;
    regs_read_arr(11)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(1).txprbssel;
    regs_read_arr(14)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(1);
    regs_read_arr(14)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(1);
    regs_read_arr(14)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(1);
    regs_read_arr(14)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(1);
    regs_read_arr(14)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(1).powergood;
    regs_read_arr(14)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(1).cplllock;
    regs_read_arr(14)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(1).cpllrefclklost;
    regs_read_arr(15)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(1);
    regs_read_arr(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(2);
    regs_read_arr(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(2);
    regs_read_arr(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(2).txpolarity;
    regs_read_arr(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(2).rxpolarity;
    regs_read_arr(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_LOOPBACK_BIT) <= loopback_arr(2);
    regs_read_arr(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(2).txinhibit;
    regs_read_arr(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(2).rxlpmen;
    regs_read_arr(18)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(2).txdiffctrl;
    regs_read_arr(18)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(2).txprecursor;
    regs_read_arr(18)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(2).txpostcursor;
    regs_read_arr(18)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(2).txmaincursor;
    regs_read_arr(19)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(2).rxprbssel;
    regs_read_arr(19)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(2).txprbssel;
    regs_read_arr(22)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(2);
    regs_read_arr(22)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(2);
    regs_read_arr(22)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(2);
    regs_read_arr(22)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(2);
    regs_read_arr(22)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(2).powergood;
    regs_read_arr(22)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(2).cplllock;
    regs_read_arr(22)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(2).cpllrefclklost;
    regs_read_arr(23)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(2);
    regs_read_arr(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(3);
    regs_read_arr(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(3);
    regs_read_arr(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(3).txpolarity;
    regs_read_arr(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(3).rxpolarity;
    regs_read_arr(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_LOOPBACK_BIT) <= loopback_arr(3);
    regs_read_arr(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(3).txinhibit;
    regs_read_arr(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(3).rxlpmen;
    regs_read_arr(26)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(3).txdiffctrl;
    regs_read_arr(26)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(3).txprecursor;
    regs_read_arr(26)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(3).txpostcursor;
    regs_read_arr(26)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(3).txmaincursor;
    regs_read_arr(27)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(3).rxprbssel;
    regs_read_arr(27)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(3).txprbssel;
    regs_read_arr(30)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(3);
    regs_read_arr(30)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(3);
    regs_read_arr(30)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(3);
    regs_read_arr(30)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(3);
    regs_read_arr(30)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(3).powergood;
    regs_read_arr(30)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(3).cplllock;
    regs_read_arr(30)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(3).cpllrefclklost;
    regs_read_arr(31)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(3);
    regs_read_arr(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(4);
    regs_read_arr(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(4);
    regs_read_arr(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(4).txpolarity;
    regs_read_arr(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(4).rxpolarity;
    regs_read_arr(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_LOOPBACK_BIT) <= loopback_arr(4);
    regs_read_arr(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(4).txinhibit;
    regs_read_arr(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(4).rxlpmen;
    regs_read_arr(34)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(4).txdiffctrl;
    regs_read_arr(34)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(4).txprecursor;
    regs_read_arr(34)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(4).txpostcursor;
    regs_read_arr(34)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(4).txmaincursor;
    regs_read_arr(35)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(4).rxprbssel;
    regs_read_arr(35)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(4).txprbssel;
    regs_read_arr(38)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(4);
    regs_read_arr(38)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(4);
    regs_read_arr(38)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(4);
    regs_read_arr(38)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(4);
    regs_read_arr(38)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(4).powergood;
    regs_read_arr(38)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(4).cplllock;
    regs_read_arr(38)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(4).cpllrefclklost;
    regs_read_arr(39)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(4);
    regs_read_arr(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(5);
    regs_read_arr(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(5);
    regs_read_arr(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(5).txpolarity;
    regs_read_arr(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(5).rxpolarity;
    regs_read_arr(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_LOOPBACK_BIT) <= loopback_arr(5);
    regs_read_arr(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(5).txinhibit;
    regs_read_arr(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(5).rxlpmen;
    regs_read_arr(42)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(5).txdiffctrl;
    regs_read_arr(42)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(5).txprecursor;
    regs_read_arr(42)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(5).txpostcursor;
    regs_read_arr(42)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(5).txmaincursor;
    regs_read_arr(43)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(5).rxprbssel;
    regs_read_arr(43)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(5).txprbssel;
    regs_read_arr(46)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(5);
    regs_read_arr(46)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(5);
    regs_read_arr(46)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(5);
    regs_read_arr(46)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(5);
    regs_read_arr(46)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(5).powergood;
    regs_read_arr(46)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(5).cplllock;
    regs_read_arr(46)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(5).cpllrefclklost;
    regs_read_arr(47)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(5);
    regs_read_arr(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(6);
    regs_read_arr(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(6);
    regs_read_arr(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(6).txpolarity;
    regs_read_arr(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(6).rxpolarity;
    regs_read_arr(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_LOOPBACK_BIT) <= loopback_arr(6);
    regs_read_arr(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(6).txinhibit;
    regs_read_arr(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(6).rxlpmen;
    regs_read_arr(50)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(6).txdiffctrl;
    regs_read_arr(50)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(6).txprecursor;
    regs_read_arr(50)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(6).txpostcursor;
    regs_read_arr(50)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(6).txmaincursor;
    regs_read_arr(51)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(6).rxprbssel;
    regs_read_arr(51)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(6).txprbssel;
    regs_read_arr(54)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(6);
    regs_read_arr(54)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(6);
    regs_read_arr(54)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(6);
    regs_read_arr(54)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(6);
    regs_read_arr(54)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(6).powergood;
    regs_read_arr(54)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(6).cplllock;
    regs_read_arr(54)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(6).cpllrefclklost;
    regs_read_arr(55)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(6);
    regs_read_arr(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(7);
    regs_read_arr(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(7);
    regs_read_arr(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(7).txpolarity;
    regs_read_arr(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(7).rxpolarity;
    regs_read_arr(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_LOOPBACK_BIT) <= loopback_arr(7);
    regs_read_arr(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(7).txinhibit;
    regs_read_arr(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(7).rxlpmen;
    regs_read_arr(58)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(7).txdiffctrl;
    regs_read_arr(58)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(7).txprecursor;
    regs_read_arr(58)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(7).txpostcursor;
    regs_read_arr(58)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(7).txmaincursor;
    regs_read_arr(59)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(7).rxprbssel;
    regs_read_arr(59)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(7).txprbssel;
    regs_read_arr(62)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(7);
    regs_read_arr(62)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(7);
    regs_read_arr(62)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(7);
    regs_read_arr(62)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(7);
    regs_read_arr(62)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(7).powergood;
    regs_read_arr(62)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(7).cplllock;
    regs_read_arr(62)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(7).cpllrefclklost;
    regs_read_arr(63)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(7);
    regs_read_arr(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(8);
    regs_read_arr(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(8);
    regs_read_arr(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(8).txpolarity;
    regs_read_arr(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(8).rxpolarity;
    regs_read_arr(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_LOOPBACK_BIT) <= loopback_arr(8);
    regs_read_arr(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(8).txinhibit;
    regs_read_arr(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(8).rxlpmen;
    regs_read_arr(66)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(8).txdiffctrl;
    regs_read_arr(66)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(8).txprecursor;
    regs_read_arr(66)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(8).txpostcursor;
    regs_read_arr(66)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(8).txmaincursor;
    regs_read_arr(67)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(8).rxprbssel;
    regs_read_arr(67)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(8).txprbssel;
    regs_read_arr(70)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(8);
    regs_read_arr(70)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(8);
    regs_read_arr(70)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(8);
    regs_read_arr(70)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(8);
    regs_read_arr(70)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(8).powergood;
    regs_read_arr(70)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(8).cplllock;
    regs_read_arr(70)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(8).cpllrefclklost;
    regs_read_arr(71)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(8);
    regs_read_arr(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(9);
    regs_read_arr(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(9);
    regs_read_arr(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(9).txpolarity;
    regs_read_arr(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(9).rxpolarity;
    regs_read_arr(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_LOOPBACK_BIT) <= loopback_arr(9);
    regs_read_arr(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(9).txinhibit;
    regs_read_arr(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(9).rxlpmen;
    regs_read_arr(74)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(9).txdiffctrl;
    regs_read_arr(74)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(9).txprecursor;
    regs_read_arr(74)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(9).txpostcursor;
    regs_read_arr(74)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(9).txmaincursor;
    regs_read_arr(75)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(9).rxprbssel;
    regs_read_arr(75)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(9).txprbssel;
    regs_read_arr(78)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(9);
    regs_read_arr(78)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(9);
    regs_read_arr(78)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(9);
    regs_read_arr(78)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(9);
    regs_read_arr(78)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(9).powergood;
    regs_read_arr(78)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(9).cplllock;
    regs_read_arr(78)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(9).cpllrefclklost;
    regs_read_arr(79)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(9);
    regs_read_arr(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(10);
    regs_read_arr(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(10);
    regs_read_arr(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(10).txpolarity;
    regs_read_arr(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(10).rxpolarity;
    regs_read_arr(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_LOOPBACK_BIT) <= loopback_arr(10);
    regs_read_arr(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(10).txinhibit;
    regs_read_arr(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(10).rxlpmen;
    regs_read_arr(82)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(10).txdiffctrl;
    regs_read_arr(82)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(10).txprecursor;
    regs_read_arr(82)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(10).txpostcursor;
    regs_read_arr(82)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(10).txmaincursor;
    regs_read_arr(83)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(10).rxprbssel;
    regs_read_arr(83)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(10).txprbssel;
    regs_read_arr(86)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(10);
    regs_read_arr(86)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(10);
    regs_read_arr(86)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(10);
    regs_read_arr(86)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(10);
    regs_read_arr(86)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(10).powergood;
    regs_read_arr(86)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(10).cplllock;
    regs_read_arr(86)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(10).cpllrefclklost;
    regs_read_arr(87)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(10);
    regs_read_arr(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(11);
    regs_read_arr(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(11);
    regs_read_arr(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(11).txpolarity;
    regs_read_arr(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(11).rxpolarity;
    regs_read_arr(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_LOOPBACK_BIT) <= loopback_arr(11);
    regs_read_arr(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(11).txinhibit;
    regs_read_arr(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(11).rxlpmen;
    regs_read_arr(90)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(11).txdiffctrl;
    regs_read_arr(90)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(11).txprecursor;
    regs_read_arr(90)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(11).txpostcursor;
    regs_read_arr(90)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(11).txmaincursor;
    regs_read_arr(91)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(11).rxprbssel;
    regs_read_arr(91)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(11).txprbssel;
    regs_read_arr(94)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(11);
    regs_read_arr(94)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(11);
    regs_read_arr(94)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(11);
    regs_read_arr(94)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(11);
    regs_read_arr(94)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(11).powergood;
    regs_read_arr(94)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(11).cplllock;
    regs_read_arr(94)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(11).cpllrefclklost;
    regs_read_arr(95)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(11);
    regs_read_arr(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(12);
    regs_read_arr(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(12);
    regs_read_arr(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(12).txpolarity;
    regs_read_arr(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(12).rxpolarity;
    regs_read_arr(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_LOOPBACK_BIT) <= loopback_arr(12);
    regs_read_arr(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(12).txinhibit;
    regs_read_arr(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(12).rxlpmen;
    regs_read_arr(98)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(12).txdiffctrl;
    regs_read_arr(98)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(12).txprecursor;
    regs_read_arr(98)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(12).txpostcursor;
    regs_read_arr(98)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(12).txmaincursor;
    regs_read_arr(99)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(12).rxprbssel;
    regs_read_arr(99)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(12).txprbssel;
    regs_read_arr(102)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(12);
    regs_read_arr(102)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(12);
    regs_read_arr(102)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(12);
    regs_read_arr(102)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(12);
    regs_read_arr(102)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(12).powergood;
    regs_read_arr(102)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(12).cplllock;
    regs_read_arr(102)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(12).cpllrefclklost;
    regs_read_arr(103)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(12);
    regs_read_arr(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(13);
    regs_read_arr(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(13);
    regs_read_arr(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(13).txpolarity;
    regs_read_arr(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(13).rxpolarity;
    regs_read_arr(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_LOOPBACK_BIT) <= loopback_arr(13);
    regs_read_arr(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(13).txinhibit;
    regs_read_arr(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(13).rxlpmen;
    regs_read_arr(106)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(13).txdiffctrl;
    regs_read_arr(106)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(13).txprecursor;
    regs_read_arr(106)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(13).txpostcursor;
    regs_read_arr(106)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(13).txmaincursor;
    regs_read_arr(107)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(13).rxprbssel;
    regs_read_arr(107)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(13).txprbssel;
    regs_read_arr(110)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(13);
    regs_read_arr(110)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(13);
    regs_read_arr(110)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(13);
    regs_read_arr(110)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(13);
    regs_read_arr(110)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(13).powergood;
    regs_read_arr(110)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(13).cplllock;
    regs_read_arr(110)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(13).cpllrefclklost;
    regs_read_arr(111)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(13);
    regs_read_arr(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(14);
    regs_read_arr(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(14);
    regs_read_arr(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(14).txpolarity;
    regs_read_arr(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(14).rxpolarity;
    regs_read_arr(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_LOOPBACK_BIT) <= loopback_arr(14);
    regs_read_arr(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(14).txinhibit;
    regs_read_arr(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(14).rxlpmen;
    regs_read_arr(114)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(14).txdiffctrl;
    regs_read_arr(114)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(14).txprecursor;
    regs_read_arr(114)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(14).txpostcursor;
    regs_read_arr(114)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(14).txmaincursor;
    regs_read_arr(115)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(14).rxprbssel;
    regs_read_arr(115)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(14).txprbssel;
    regs_read_arr(118)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(14);
    regs_read_arr(118)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(14);
    regs_read_arr(118)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(14);
    regs_read_arr(118)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(14);
    regs_read_arr(118)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(14).powergood;
    regs_read_arr(118)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(14).cplllock;
    regs_read_arr(118)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(14).cpllrefclklost;
    regs_read_arr(119)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(14);
    regs_read_arr(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_POWERDOWN_BIT) <= txpd_arr(15);
    regs_read_arr(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_POWERDOWN_BIT) <= rxpd_arr(15);
    regs_read_arr(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_POLARITY_BIT) <= tx_slow_ctrl_arr(15).txpolarity;
    regs_read_arr(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_POLARITY_BIT) <= rx_slow_ctrl_arr(15).rxpolarity;
    regs_read_arr(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_LOOPBACK_BIT) <= loopback_arr(15);
    regs_read_arr(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_INHIBIT_BIT) <= tx_slow_ctrl_arr(15).txinhibit;
    regs_read_arr(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_LOW_POWER_MODE_BIT) <= rx_slow_ctrl_arr(15).rxlpmen;
    regs_read_arr(122)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_DIFF_CTRL_LSB) <= tx_slow_ctrl_arr(15).txdiffctrl;
    regs_read_arr(122)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_PRE_CURSOR_LSB) <= tx_slow_ctrl_arr(15).txprecursor;
    regs_read_arr(122)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_POST_CURSOR_LSB) <= tx_slow_ctrl_arr(15).txpostcursor;
    regs_read_arr(122)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_MAIN_CURSOR_LSB) <= tx_slow_ctrl_arr(15).txmaincursor;
    regs_read_arr(123)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_PRBS_SEL_LSB) <= rx_slow_ctrl_arr(15).rxprbssel;
    regs_read_arr(123)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_PRBS_SEL_LSB) <= tx_slow_ctrl_arr(15).txprbssel;
    regs_read_arr(126)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_STATUS_TX_RESET_DONE_BIT) <= tx_reset_done_arr_i(15);
    regs_read_arr(126)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_STATUS_RX_RESET_DONE_BIT) <= rx_reset_done_arr_i(15);
    regs_read_arr(126)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_STATUS_TX_PHALIGN_DONE_BIT) <= tx_phalign_done_arr_i(15);
    regs_read_arr(126)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_STATUS_RX_PHALIGN_DONE_BIT) <= rx_phalign_done_arr_i(15);
    regs_read_arr(126)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_STATUS_POWER_GOOD_BIT) <= misc_status_arr_i(15).powergood;
    regs_read_arr(126)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_STATUS_CPLL_LOCKED_BIT) <= cpll_status_arr_i(15).cplllock;
    regs_read_arr(126)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_STATUS_CPLL_REF_CLK_LOST_BIT) <= cpll_status_arr_i(15).cpllrefclklost;
    regs_read_arr(127)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_STATUS_PRBS_ERROR_CNT_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_STATUS_PRBS_ERROR_CNT_LSB) <= prbs_err_cnt_sync_arr(15);

    -- Connect write signals
    txpd_arr(0) <= regs_write_arr(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(0) <= regs_write_arr(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(0).txpolarity <= regs_write_arr(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(0).rxpolarity <= regs_write_arr(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_POLARITY_BIT);
    loopback_arr(0) <= regs_write_arr(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(0).txinhibit <= regs_write_arr(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(0).rxlpmen <= regs_write_arr(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(0).txdiffctrl <= regs_write_arr(2)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(0).txprecursor <= regs_write_arr(2)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(0).txpostcursor <= regs_write_arr(2)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(0).txmaincursor <= regs_write_arr(2)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(0).rxprbssel <= regs_write_arr(3)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(0).txprbssel <= regs_write_arr(3)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_PRBS_SEL_LSB);
    txpd_arr(1) <= regs_write_arr(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(1) <= regs_write_arr(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(1).txpolarity <= regs_write_arr(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(1).rxpolarity <= regs_write_arr(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_POLARITY_BIT);
    loopback_arr(1) <= regs_write_arr(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(1).txinhibit <= regs_write_arr(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(1).rxlpmen <= regs_write_arr(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(1).txdiffctrl <= regs_write_arr(10)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(1).txprecursor <= regs_write_arr(10)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(1).txpostcursor <= regs_write_arr(10)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(1).txmaincursor <= regs_write_arr(10)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(1).rxprbssel <= regs_write_arr(11)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(1).txprbssel <= regs_write_arr(11)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_PRBS_SEL_LSB);
    txpd_arr(2) <= regs_write_arr(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(2) <= regs_write_arr(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(2).txpolarity <= regs_write_arr(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(2).rxpolarity <= regs_write_arr(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_POLARITY_BIT);
    loopback_arr(2) <= regs_write_arr(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(2).txinhibit <= regs_write_arr(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(2).rxlpmen <= regs_write_arr(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(2).txdiffctrl <= regs_write_arr(18)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(2).txprecursor <= regs_write_arr(18)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(2).txpostcursor <= regs_write_arr(18)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(2).txmaincursor <= regs_write_arr(18)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(2).rxprbssel <= regs_write_arr(19)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(2).txprbssel <= regs_write_arr(19)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_PRBS_SEL_LSB);
    txpd_arr(3) <= regs_write_arr(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(3) <= regs_write_arr(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(3).txpolarity <= regs_write_arr(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(3).rxpolarity <= regs_write_arr(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_POLARITY_BIT);
    loopback_arr(3) <= regs_write_arr(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(3).txinhibit <= regs_write_arr(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(3).rxlpmen <= regs_write_arr(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(3).txdiffctrl <= regs_write_arr(26)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(3).txprecursor <= regs_write_arr(26)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(3).txpostcursor <= regs_write_arr(26)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(3).txmaincursor <= regs_write_arr(26)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(3).rxprbssel <= regs_write_arr(27)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(3).txprbssel <= regs_write_arr(27)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_PRBS_SEL_LSB);
    txpd_arr(4) <= regs_write_arr(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(4) <= regs_write_arr(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(4).txpolarity <= regs_write_arr(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(4).rxpolarity <= regs_write_arr(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_POLARITY_BIT);
    loopback_arr(4) <= regs_write_arr(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(4).txinhibit <= regs_write_arr(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(4).rxlpmen <= regs_write_arr(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(4).txdiffctrl <= regs_write_arr(34)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(4).txprecursor <= regs_write_arr(34)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(4).txpostcursor <= regs_write_arr(34)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(4).txmaincursor <= regs_write_arr(34)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(4).rxprbssel <= regs_write_arr(35)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(4).txprbssel <= regs_write_arr(35)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_PRBS_SEL_LSB);
    txpd_arr(5) <= regs_write_arr(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(5) <= regs_write_arr(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(5).txpolarity <= regs_write_arr(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(5).rxpolarity <= regs_write_arr(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_POLARITY_BIT);
    loopback_arr(5) <= regs_write_arr(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(5).txinhibit <= regs_write_arr(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(5).rxlpmen <= regs_write_arr(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(5).txdiffctrl <= regs_write_arr(42)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(5).txprecursor <= regs_write_arr(42)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(5).txpostcursor <= regs_write_arr(42)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(5).txmaincursor <= regs_write_arr(42)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(5).rxprbssel <= regs_write_arr(43)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(5).txprbssel <= regs_write_arr(43)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_PRBS_SEL_LSB);
    txpd_arr(6) <= regs_write_arr(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(6) <= regs_write_arr(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(6).txpolarity <= regs_write_arr(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(6).rxpolarity <= regs_write_arr(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_POLARITY_BIT);
    loopback_arr(6) <= regs_write_arr(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(6).txinhibit <= regs_write_arr(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(6).rxlpmen <= regs_write_arr(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(6).txdiffctrl <= regs_write_arr(50)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(6).txprecursor <= regs_write_arr(50)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(6).txpostcursor <= regs_write_arr(50)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(6).txmaincursor <= regs_write_arr(50)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(6).rxprbssel <= regs_write_arr(51)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(6).txprbssel <= regs_write_arr(51)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_PRBS_SEL_LSB);
    txpd_arr(7) <= regs_write_arr(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(7) <= regs_write_arr(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(7).txpolarity <= regs_write_arr(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(7).rxpolarity <= regs_write_arr(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_POLARITY_BIT);
    loopback_arr(7) <= regs_write_arr(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(7).txinhibit <= regs_write_arr(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(7).rxlpmen <= regs_write_arr(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(7).txdiffctrl <= regs_write_arr(58)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(7).txprecursor <= regs_write_arr(58)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(7).txpostcursor <= regs_write_arr(58)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(7).txmaincursor <= regs_write_arr(58)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(7).rxprbssel <= regs_write_arr(59)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(7).txprbssel <= regs_write_arr(59)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_PRBS_SEL_LSB);
    txpd_arr(8) <= regs_write_arr(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(8) <= regs_write_arr(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(8).txpolarity <= regs_write_arr(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(8).rxpolarity <= regs_write_arr(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_POLARITY_BIT);
    loopback_arr(8) <= regs_write_arr(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(8).txinhibit <= regs_write_arr(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(8).rxlpmen <= regs_write_arr(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(8).txdiffctrl <= regs_write_arr(66)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(8).txprecursor <= regs_write_arr(66)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(8).txpostcursor <= regs_write_arr(66)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(8).txmaincursor <= regs_write_arr(66)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(8).rxprbssel <= regs_write_arr(67)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(8).txprbssel <= regs_write_arr(67)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_PRBS_SEL_LSB);
    txpd_arr(9) <= regs_write_arr(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(9) <= regs_write_arr(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(9).txpolarity <= regs_write_arr(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(9).rxpolarity <= regs_write_arr(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_POLARITY_BIT);
    loopback_arr(9) <= regs_write_arr(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(9).txinhibit <= regs_write_arr(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(9).rxlpmen <= regs_write_arr(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(9).txdiffctrl <= regs_write_arr(74)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(9).txprecursor <= regs_write_arr(74)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(9).txpostcursor <= regs_write_arr(74)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(9).txmaincursor <= regs_write_arr(74)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(9).rxprbssel <= regs_write_arr(75)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(9).txprbssel <= regs_write_arr(75)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_PRBS_SEL_LSB);
    txpd_arr(10) <= regs_write_arr(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(10) <= regs_write_arr(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(10).txpolarity <= regs_write_arr(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(10).rxpolarity <= regs_write_arr(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_POLARITY_BIT);
    loopback_arr(10) <= regs_write_arr(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(10).txinhibit <= regs_write_arr(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(10).rxlpmen <= regs_write_arr(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(10).txdiffctrl <= regs_write_arr(82)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(10).txprecursor <= regs_write_arr(82)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(10).txpostcursor <= regs_write_arr(82)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(10).txmaincursor <= regs_write_arr(82)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(10).rxprbssel <= regs_write_arr(83)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(10).txprbssel <= regs_write_arr(83)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_PRBS_SEL_LSB);
    txpd_arr(11) <= regs_write_arr(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(11) <= regs_write_arr(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(11).txpolarity <= regs_write_arr(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(11).rxpolarity <= regs_write_arr(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_POLARITY_BIT);
    loopback_arr(11) <= regs_write_arr(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(11).txinhibit <= regs_write_arr(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(11).rxlpmen <= regs_write_arr(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(11).txdiffctrl <= regs_write_arr(90)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(11).txprecursor <= regs_write_arr(90)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(11).txpostcursor <= regs_write_arr(90)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(11).txmaincursor <= regs_write_arr(90)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(11).rxprbssel <= regs_write_arr(91)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(11).txprbssel <= regs_write_arr(91)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_PRBS_SEL_LSB);
    txpd_arr(12) <= regs_write_arr(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(12) <= regs_write_arr(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(12).txpolarity <= regs_write_arr(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(12).rxpolarity <= regs_write_arr(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_POLARITY_BIT);
    loopback_arr(12) <= regs_write_arr(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(12).txinhibit <= regs_write_arr(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(12).rxlpmen <= regs_write_arr(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(12).txdiffctrl <= regs_write_arr(98)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(12).txprecursor <= regs_write_arr(98)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(12).txpostcursor <= regs_write_arr(98)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(12).txmaincursor <= regs_write_arr(98)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(12).rxprbssel <= regs_write_arr(99)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(12).txprbssel <= regs_write_arr(99)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_PRBS_SEL_LSB);
    txpd_arr(13) <= regs_write_arr(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(13) <= regs_write_arr(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(13).txpolarity <= regs_write_arr(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(13).rxpolarity <= regs_write_arr(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_POLARITY_BIT);
    loopback_arr(13) <= regs_write_arr(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(13).txinhibit <= regs_write_arr(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(13).rxlpmen <= regs_write_arr(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(13).txdiffctrl <= regs_write_arr(106)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(13).txprecursor <= regs_write_arr(106)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(13).txpostcursor <= regs_write_arr(106)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(13).txmaincursor <= regs_write_arr(106)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(13).rxprbssel <= regs_write_arr(107)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(13).txprbssel <= regs_write_arr(107)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_PRBS_SEL_LSB);
    txpd_arr(14) <= regs_write_arr(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(14) <= regs_write_arr(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(14).txpolarity <= regs_write_arr(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(14).rxpolarity <= regs_write_arr(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_POLARITY_BIT);
    loopback_arr(14) <= regs_write_arr(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(14).txinhibit <= regs_write_arr(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(14).rxlpmen <= regs_write_arr(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(14).txdiffctrl <= regs_write_arr(114)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(14).txprecursor <= regs_write_arr(114)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(14).txpostcursor <= regs_write_arr(114)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(14).txmaincursor <= regs_write_arr(114)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(14).rxprbssel <= regs_write_arr(115)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(14).txprbssel <= regs_write_arr(115)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_PRBS_SEL_LSB);
    txpd_arr(15) <= regs_write_arr(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_POWERDOWN_BIT);
    rxpd_arr(15) <= regs_write_arr(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_POWERDOWN_BIT);
    tx_slow_ctrl_arr(15).txpolarity <= regs_write_arr(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_POLARITY_BIT);
    rx_slow_ctrl_arr(15).rxpolarity <= regs_write_arr(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_POLARITY_BIT);
    loopback_arr(15) <= regs_write_arr(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_LOOPBACK_BIT);
    tx_slow_ctrl_arr(15).txinhibit <= regs_write_arr(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_INHIBIT_BIT);
    rx_slow_ctrl_arr(15).rxlpmen <= regs_write_arr(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_LOW_POWER_MODE_BIT);
    tx_slow_ctrl_arr(15).txdiffctrl <= regs_write_arr(122)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_DIFF_CTRL_LSB);
    tx_slow_ctrl_arr(15).txprecursor <= regs_write_arr(122)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_PRE_CURSOR_LSB);
    tx_slow_ctrl_arr(15).txpostcursor <= regs_write_arr(122)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_POST_CURSOR_LSB);
    tx_slow_ctrl_arr(15).txmaincursor <= regs_write_arr(122)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_MAIN_CURSOR_LSB);
    rx_slow_ctrl_arr(15).rxprbssel <= regs_write_arr(123)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_PRBS_SEL_LSB);
    tx_slow_ctrl_arr(15).txprbssel <= regs_write_arr(123)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_PRBS_SEL_LSB);

    -- Connect write pulse signals
    reset_arr(0) <= regs_write_pulse_arr(0);
    tx_slow_ctrl_arr(0).txprbsforceerr <= regs_write_pulse_arr(4);
    prbs_err_reset_arr(0) <= regs_write_pulse_arr(5);
    reset_arr(1) <= regs_write_pulse_arr(8);
    tx_slow_ctrl_arr(1).txprbsforceerr <= regs_write_pulse_arr(12);
    prbs_err_reset_arr(1) <= regs_write_pulse_arr(13);
    reset_arr(2) <= regs_write_pulse_arr(16);
    tx_slow_ctrl_arr(2).txprbsforceerr <= regs_write_pulse_arr(20);
    prbs_err_reset_arr(2) <= regs_write_pulse_arr(21);
    reset_arr(3) <= regs_write_pulse_arr(24);
    tx_slow_ctrl_arr(3).txprbsforceerr <= regs_write_pulse_arr(28);
    prbs_err_reset_arr(3) <= regs_write_pulse_arr(29);
    reset_arr(4) <= regs_write_pulse_arr(32);
    tx_slow_ctrl_arr(4).txprbsforceerr <= regs_write_pulse_arr(36);
    prbs_err_reset_arr(4) <= regs_write_pulse_arr(37);
    reset_arr(5) <= regs_write_pulse_arr(40);
    tx_slow_ctrl_arr(5).txprbsforceerr <= regs_write_pulse_arr(44);
    prbs_err_reset_arr(5) <= regs_write_pulse_arr(45);
    reset_arr(6) <= regs_write_pulse_arr(48);
    tx_slow_ctrl_arr(6).txprbsforceerr <= regs_write_pulse_arr(52);
    prbs_err_reset_arr(6) <= regs_write_pulse_arr(53);
    reset_arr(7) <= regs_write_pulse_arr(56);
    tx_slow_ctrl_arr(7).txprbsforceerr <= regs_write_pulse_arr(60);
    prbs_err_reset_arr(7) <= regs_write_pulse_arr(61);
    reset_arr(8) <= regs_write_pulse_arr(64);
    tx_slow_ctrl_arr(8).txprbsforceerr <= regs_write_pulse_arr(68);
    prbs_err_reset_arr(8) <= regs_write_pulse_arr(69);
    reset_arr(9) <= regs_write_pulse_arr(72);
    tx_slow_ctrl_arr(9).txprbsforceerr <= regs_write_pulse_arr(76);
    prbs_err_reset_arr(9) <= regs_write_pulse_arr(77);
    reset_arr(10) <= regs_write_pulse_arr(80);
    tx_slow_ctrl_arr(10).txprbsforceerr <= regs_write_pulse_arr(84);
    prbs_err_reset_arr(10) <= regs_write_pulse_arr(85);
    reset_arr(11) <= regs_write_pulse_arr(88);
    tx_slow_ctrl_arr(11).txprbsforceerr <= regs_write_pulse_arr(92);
    prbs_err_reset_arr(11) <= regs_write_pulse_arr(93);
    reset_arr(12) <= regs_write_pulse_arr(96);
    tx_slow_ctrl_arr(12).txprbsforceerr <= regs_write_pulse_arr(100);
    prbs_err_reset_arr(12) <= regs_write_pulse_arr(101);
    reset_arr(13) <= regs_write_pulse_arr(104);
    tx_slow_ctrl_arr(13).txprbsforceerr <= regs_write_pulse_arr(108);
    prbs_err_reset_arr(13) <= regs_write_pulse_arr(109);
    reset_arr(14) <= regs_write_pulse_arr(112);
    tx_slow_ctrl_arr(14).txprbsforceerr <= regs_write_pulse_arr(116);
    prbs_err_reset_arr(14) <= regs_write_pulse_arr(117);
    reset_arr(15) <= regs_write_pulse_arr(120);
    tx_slow_ctrl_arr(15).txprbsforceerr <= regs_write_pulse_arr(124);
    prbs_err_reset_arr(15) <= regs_write_pulse_arr(125);

    -- Connect write done signals

    -- Connect read pulse signals

    -- Connect read ready signals

    -- Defaults
    regs_defaults(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(1)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(2)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(2)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(2)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(2)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(3)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(3)(REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_0_CTRL_TX_PRBS_SEL_DEFAULT;
    regs_defaults(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(9)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(10)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(10)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(10)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(10)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(11)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(11)(REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_1_CTRL_TX_PRBS_SEL_DEFAULT;
    regs_defaults(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(17)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(18)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(18)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(18)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(18)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(19)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(19)(REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_2_CTRL_TX_PRBS_SEL_DEFAULT;
    regs_defaults(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(25)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(26)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(26)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(26)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(26)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(27)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(27)(REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_3_CTRL_TX_PRBS_SEL_DEFAULT;
    regs_defaults(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(33)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(34)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(34)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(34)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(34)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(35)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(35)(REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_4_CTRL_TX_PRBS_SEL_DEFAULT;
    regs_defaults(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(41)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(42)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(42)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(42)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(42)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(43)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(43)(REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_5_CTRL_TX_PRBS_SEL_DEFAULT;
    regs_defaults(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(49)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(50)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(50)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(50)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(50)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(51)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(51)(REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_6_CTRL_TX_PRBS_SEL_DEFAULT;
    regs_defaults(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(57)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(58)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(58)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(58)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(58)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(59)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(59)(REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_7_CTRL_TX_PRBS_SEL_DEFAULT;
    regs_defaults(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(65)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(66)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(66)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(66)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(66)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(67)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(67)(REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_8_CTRL_TX_PRBS_SEL_DEFAULT;
    regs_defaults(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(73)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(74)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(74)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(74)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(74)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(75)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(75)(REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_9_CTRL_TX_PRBS_SEL_DEFAULT;
    regs_defaults(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(81)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(82)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(82)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(82)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(82)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(83)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(83)(REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_10_CTRL_TX_PRBS_SEL_DEFAULT;
    regs_defaults(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(89)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(90)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(90)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(90)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(90)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(91)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(91)(REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_11_CTRL_TX_PRBS_SEL_DEFAULT;
    regs_defaults(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(97)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(98)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(98)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(98)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(98)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(99)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(99)(REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_12_CTRL_TX_PRBS_SEL_DEFAULT;
    regs_defaults(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(105)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(106)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(106)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(106)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(106)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(107)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(107)(REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_13_CTRL_TX_PRBS_SEL_DEFAULT;
    regs_defaults(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(113)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(114)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(114)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(114)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(114)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(115)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(115)(REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_14_CTRL_TX_PRBS_SEL_DEFAULT;
    regs_defaults(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_POWERDOWN_DEFAULT;
    regs_defaults(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_POWERDOWN_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_POWERDOWN_DEFAULT;
    regs_defaults(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_POLARITY_DEFAULT;
    regs_defaults(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_POLARITY_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_POLARITY_DEFAULT;
    regs_defaults(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_LOOPBACK_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_LOOPBACK_DEFAULT;
    regs_defaults(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_INHIBIT_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_INHIBIT_DEFAULT;
    regs_defaults(121)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_LOW_POWER_MODE_BIT) <= REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_LOW_POWER_MODE_DEFAULT;
    regs_defaults(122)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_DIFF_CTRL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_DIFF_CTRL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_DIFF_CTRL_DEFAULT;
    regs_defaults(122)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_PRE_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_PRE_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_PRE_CURSOR_DEFAULT;
    regs_defaults(122)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_POST_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_POST_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_POST_CURSOR_DEFAULT;
    regs_defaults(122)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_MAIN_CURSOR_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_MAIN_CURSOR_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_MAIN_CURSOR_DEFAULT;
    regs_defaults(123)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_RX_PRBS_SEL_DEFAULT;
    regs_defaults(123)(REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_PRBS_SEL_MSB downto REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_PRBS_SEL_LSB) <= REG_OPTICAL_LINKS_MGT_CHANNEL_15_CTRL_TX_PRBS_SEL_DEFAULT;

    -- Define writable regs
    regs_writable_arr(1) <= '1';
    regs_writable_arr(2) <= '1';
    regs_writable_arr(3) <= '1';
    regs_writable_arr(9) <= '1';
    regs_writable_arr(10) <= '1';
    regs_writable_arr(11) <= '1';
    regs_writable_arr(17) <= '1';
    regs_writable_arr(18) <= '1';
    regs_writable_arr(19) <= '1';
    regs_writable_arr(25) <= '1';
    regs_writable_arr(26) <= '1';
    regs_writable_arr(27) <= '1';
    regs_writable_arr(33) <= '1';
    regs_writable_arr(34) <= '1';
    regs_writable_arr(35) <= '1';
    regs_writable_arr(41) <= '1';
    regs_writable_arr(42) <= '1';
    regs_writable_arr(43) <= '1';
    regs_writable_arr(49) <= '1';
    regs_writable_arr(50) <= '1';
    regs_writable_arr(51) <= '1';
    regs_writable_arr(57) <= '1';
    regs_writable_arr(58) <= '1';
    regs_writable_arr(59) <= '1';
    regs_writable_arr(65) <= '1';
    regs_writable_arr(66) <= '1';
    regs_writable_arr(67) <= '1';
    regs_writable_arr(73) <= '1';
    regs_writable_arr(74) <= '1';
    regs_writable_arr(75) <= '1';
    regs_writable_arr(81) <= '1';
    regs_writable_arr(82) <= '1';
    regs_writable_arr(83) <= '1';
    regs_writable_arr(89) <= '1';
    regs_writable_arr(90) <= '1';
    regs_writable_arr(91) <= '1';
    regs_writable_arr(97) <= '1';
    regs_writable_arr(98) <= '1';
    regs_writable_arr(99) <= '1';
    regs_writable_arr(105) <= '1';
    regs_writable_arr(106) <= '1';
    regs_writable_arr(107) <= '1';
    regs_writable_arr(113) <= '1';
    regs_writable_arr(114) <= '1';
    regs_writable_arr(115) <= '1';
    regs_writable_arr(121) <= '1';
    regs_writable_arr(122) <= '1';
    regs_writable_arr(123) <= '1';

    --==== Registers end ============================================================================

end mgt_slow_control_arch;
