library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package tmr_pkg is
  constant EN_TMR : integer := 1;
end tmr_pkg;
