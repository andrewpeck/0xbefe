------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    15:04 2016-05-10
-- Module Name:    GEM System Registers
-- Description:    this module provides registers for GEM system-wide setting  
------------------------------------------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_misc.all;

use work.ipbus.all;
use work.common_pkg.all;
use work.gem_pkg.all;
use work.registers.all;
use work.ttc_pkg.all;
use work.gem_board_config_package.all;

entity gem_system_regs is
generic(
    g_NUM_IPB_MON_SLAVES     : integer;
    
    -- Firmware version, date, time, git sha
    g_FW_DATE            : std_logic_vector (31 downto 0);
    g_FW_TIME            : std_logic_vector (31 downto 0);
    g_FW_VER             : std_logic_vector (31 downto 0);
    g_FW_SHA             : std_logic_vector (31 downto 0);
    
    --remove later
    g_NUM_OF_OHs                : integer            
);
port(
    
    reset_i                     : in std_logic;

    ttc_clks_i                  : in t_ttc_clks;

    ipb_clk_i                   : in std_logic;
    ipb_reset_i                 : in std_logic;
    
    ipb_mosi_i                  : in ipb_wbus;
    ipb_miso_o                  : out ipb_rbus;
    ipb_mon_miso_arr_i          : ipb_rbus_array(g_NUM_IPB_MON_SLAVES - 1 downto 0);
    
    board_id_o                  : out std_logic_vector(15 downto 0);

    loopback_gbt_test_en_o      : out std_logic;
    use_v3b_elink_mapping_o     : out std_logic;
    use_vfat_addressing_o       : out std_logic;

    vfat3_sc_only_mode_o        : out std_logic;
    manual_link_reset_o         : out std_logic;
    global_reset_o              : out std_logic;
    gbt_reset_o                 : out std_logic;
    manual_ipbus_reset_o        : out std_logic;
    
    gemloader_stats_i           : in  t_gem_loader_stats;
    gemloader_cfg_o             : out t_gem_loader_cfg;
    
    vfat3_sbits_arr_i           : in t_vfat3_sbits_arr(g_NUM_OF_OHs - 1 downto 0)
    
);
end gem_system_regs;

architecture gem_system_regs_arch of gem_system_regs is

    signal reset_cnt                : std_logic := '0';
    
    signal board_id                 : std_logic_vector(15 downto 0) := (others => '0');
    signal gem_station              : integer range 0 to 2;
    signal num_of_oh                : std_logic_vector(4 downto 0);
    signal board_type               : std_logic_vector(3 downto 0);
    
    signal loopback_gbt_test_en     : std_logic;
    
    signal vfat3_sc_only_mode       : std_logic;
    
    signal use_v3b_elink_mapping    : std_logic;
    signal use_vfat_addressing      : std_logic;

    signal global_reset_timer       : integer range 0 to 100 := 0;
    signal global_reset_trig        : std_logic;

    signal ipbus_reset_timer        : integer range 0 to 100 := 0;
    signal ipbus_reset_trig         : std_logic;

    signal ipb_mon_miso_ack_arr     : std_logic_vector(g_NUM_IPB_MON_SLAVES - 1 downto 0);
    signal ipb_mon_miso_err_arr     : std_logic_vector(g_NUM_IPB_MON_SLAVES - 1 downto 0);
    signal ipb_mon_miso_ack_or      : std_logic;
    signal ipb_mon_miso_err_or      : std_logic;
    signal ipb_mon_last_trans_err   : std_logic;
    signal ipb_mon_trans_cnt        : std_logic_vector(15 downto 0);
    signal ipb_mon_err_cnt          : std_logic_vector(14 downto 0);

    signal gemloader_fw_size        : std_logic_vector(31 downto 0);
    
    signal test_sbit_me0            : std_logic_vector(31 downto 0);
    
    signal sbit_test_reset_o            : std_logic := '0' ;
    
    signal test_sbit0xe_count_me0 : std_logic_vector(31 downto 0);
    signal vfat3_sbit0xe_test : std_logic_vector(7 downto 0);
    signal test_sbit0xs_count_me0 : std_logic_vector(31 downto 0);
    signal vfat3_sbit0xs_test : std_logic;
    signal test_sel_vfat_sbit_me0 : std_logic_vector(31 downto 0);
    signal test_sel_elink_sbit_me0 : std_logic_vector(31 downto 0);
    signal test_sel_sbit_me0 : std_logic_vector(31 downto 0);

    ------ Register signals begin (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    ------ Register signals end ----------------------------------------------
    
begin

    --=== board type and configuration parameters ===--
    board_type     <= CFG_BOARD_TYPE;
    num_of_oh      <= std_logic_vector(to_unsigned(CFG_NUM_OF_OHs, 5));
    gem_station    <= CFG_GEM_STATION;
    
    
            
    --=== Tests === --
    loopback_gbt_test_en_o <= loopback_gbt_test_en; 
    
    --=== VFAT conf === --
    vfat3_sc_only_mode_o <= vfat3_sc_only_mode;
    use_v3b_elink_mapping_o <= use_v3b_elink_mapping;
    use_vfat_addressing_o <= use_vfat_addressing;

    --=== PROMless === --
    gemloader_cfg_o.firmware_size <= gemloader_fw_size;


    --=== Global resets === --
    process (ttc_clks_i.clk_40)
    begin
        if rising_edge(ttc_clks_i.clk_40) then
            if (global_reset_trig = '1') then
                global_reset_timer <= 100;
                global_reset_o <= '0';
            else
                -- wait for 50 cycles after the trigger, and then keep the reset on for 50 cycles
                if (global_reset_timer = 0) then
                    global_reset_o <= '0';
                    global_reset_timer <= 0;
                elsif (global_reset_timer > 50) then
                    global_reset_o <= '0';
                    global_reset_timer <= global_reset_timer - 1; 
                else
                    global_reset_o <= '1';
                    global_reset_timer <= global_reset_timer - 1;
                end if;
            end if;
        end if;
    end process;

    --=== IPB reset === --
    process (ttc_clks_i.clk_40)
    begin
        if rising_edge(ttc_clks_i.clk_40) then
            if (ipbus_reset_trig = '1') then
                ipbus_reset_timer <= 100;
                manual_ipbus_reset_o <= '0';
            else
                -- wait for 50 cycles after the trigger, and then keep the reset on for 50 cycles
                if (ipbus_reset_timer = 0) then
                    manual_ipbus_reset_o <= '0';
                    ipbus_reset_timer <= 0;
                elsif (ipbus_reset_timer > 50) then
                    manual_ipbus_reset_o <= '0';
                    ipbus_reset_timer <= ipbus_reset_timer - 1; 
                else
                    manual_ipbus_reset_o <= '1';
                    ipbus_reset_timer <= ipbus_reset_timer - 1;
                end if;
            end if;
        end if;
    end process;

    --=== IPB monitor === --
    process (ipb_clk_i)
    begin
        if rising_edge(ipb_clk_i) then
            for i in 0 to g_NUM_IPB_MON_SLAVES - 1 loop
                ipb_mon_miso_ack_arr(i) <= ipb_mon_miso_arr_i(i).ipb_ack;
                ipb_mon_miso_err_arr(i) <= ipb_mon_miso_arr_i(i).ipb_err;
            end loop;
            ipb_mon_miso_ack_or <= or_reduce(ipb_mon_miso_ack_arr);
            ipb_mon_miso_err_or <= or_reduce(ipb_mon_miso_err_arr);
            
            if (ipb_mon_miso_ack_or = '1') then
                ipb_mon_last_trans_err <= ipb_mon_miso_err_or;
            end if; 
        end if;
    end process;

    i_ipb_mon_trans_cnt : entity work.counter
        generic map(
            g_COUNTER_WIDTH  => 16,
            g_ALLOW_ROLLOVER => true
        )
        port map(
            ref_clk_i => ipb_clk_i,
            reset_i   => reset_i,
            en_i      => ipb_mon_miso_ack_or,
            count_o   => ipb_mon_trans_cnt
        );

    i_ipb_mon_err_cnt : entity work.counter
        generic map(
            g_COUNTER_WIDTH  => 15,
            g_ALLOW_ROLLOVER => true
        )
        port map(
            ref_clk_i => ipb_clk_i,
            reset_i   => reset_i,
            en_i      => ipb_mon_miso_err_or,
            count_o   => ipb_mon_err_cnt
        );
     
     vfat3_sbit0xe_test <= vfat3_sbits_arr_i(0)(to_integer(unsigned(test_sel_vfat_sbit_me0)))((((to_integer(unsigned(test_sel_elink_sbit_me0 )) + 1) * 8) - 1) downto (to_integer(unsigned(test_sel_elink_sbit_me0)) * 8));
     
     me0_sbit0xe_count : entity work.counter
        generic map(
            g_COUNTER_WIDTH  => 32,
            g_ALLOW_ROLLOVER => false
        )
        port map(
            ref_clk_i => ttc_clks_i.clk_40,
            reset_i   => sbit_test_reset_o,
            en_i      => vfat3_sbit0xe_test(7) or
                         vfat3_sbit0xe_test(6) or
                         vfat3_sbit0xe_test(5) or
                         vfat3_sbit0xe_test(4) or
                         vfat3_sbit0xe_test(3) or
                         vfat3_sbit0xe_test(2) or
                         vfat3_sbit0xe_test(1) or
                         vfat3_sbit0xe_test(0),
            count_o   => test_sbit0xx_count_me0
        );   
        
     vfat3_sbit0xs_test <= vfat3_sbits_arr_i(0)(to_integer(unsigned(test_sel_vfat_sbit_me0)))(to_integer(unsigned(test_sel_sbit_me0)));
     
     me0_sbit0xs_count : entity work.counter
        generic map(
            g_COUNTER_WIDTH  => 32,
            g_ALLOW_ROLLOVER => false
        )
        port map(
            ref_clk_i => ttc_clks_i.clk_40,
            reset_i   => sbit_test_reset_o,
            en_i      => vfat3_sbit0xs_test,
            count_o   => test_sbit0xs_count_me0
        );    
     
    --===============================================================================================
    -- this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    --==== Registers end ============================================================================

end gem_system_regs_arch;
