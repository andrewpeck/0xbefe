------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    2020-07-16
-- Module Name:    PROMLESS
-- Description:    This module implements the so called gemloader module which stores the frontend firmware, and streams it to the gem logic on request.
--                 This version uses the FPGA BRAM for storing the bitfile  
------------------------------------------------------------------------------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library xpm;
use xpm.vcomponents.all;

use work.ttc_pkg.all;
use work.common_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity promless is
    generic(
        g_MAX_SIZE_BYTES    : integer; -- NOTE: must be a multiple of 32KB (kilobytes) if g_MEMORY_PRIMITIVE is set to "ultra" (using UltraRAM)
        g_MEMORY_PRIMITIVE  : string := "ultra";
        g_IPB_CLK_PERIOD_NS : integer
    );
    port (
        reset_i             : in  std_logic;
        
        to_promless_i       : in  t_to_promless;
        from_promless_o     : out t_from_promless;        
        
        -- IPbus
        ipb_reset_i         : in  std_logic;
        ipb_clk_i           : in  std_logic;
        ipb_miso_o          : out ipb_rbus;
        ipb_mosi_i          : in  ipb_wbus                
    );
end promless;

architecture promless_arch of promless is

    ----==== RAM signals ====----
    
    -- port A is used by the IPbus slave (write and read), and port B is used by the loader (read-only)
    
    constant RAM_ADDR_WIDTH   : integer := 20;
    constant RAM_READ_LATENCY : integer := 8;
    
    -- Common RAM port A signals 
    signal rama_addr                : std_logic_vector(RAM_ADDR_WIDTH - 1 downto 0) := (others => '0');
    signal rama_din                 : std_logic_vector(63 downto 0) := (others => '0');
    signal rama_we                  : std_logic_vector(7 downto 0)  := (others => '0');
    signal rama_dout                : std_logic_vector(63 downto 0);

    signal rama_write_req           : std_logic;
    signal rama_read_req            : std_logic;
    signal rama_read_ready          : std_logic;
    signal rama_read_ready_pipe     : std_logic_vector(RAM_READ_LATENCY downto 0) := (others => '0');
    signal rama_write_addr          : std_logic_vector(RAM_ADDR_WIDTH downto 0) := (others => '0');
    signal rama_read_addr           : std_logic_vector(RAM_ADDR_WIDTH downto 0) := (others => '0');
    signal rama_reset_addr          : std_logic;
    signal rama_write_data          : std_logic_vector(31 downto 0) := (others => '0');
    signal rama_read_data           : std_logic_vector(31 downto 0) := (others => '0');

    -- port B signals
    signal ramb_addr                : std_logic_vector(RAM_ADDR_WIDTH - 1 downto 0) := (others => '0');
    signal ramb_dout                : std_logic_vector(63 downto 0);
    signal ramb_byte_sel            : std_logic_vector(2 downto 0) := (others => '0');
    signal ramb_byte_sel_pipe       : t_std3_array(RAM_READ_LATENCY downto 0) := (others => (others => '0'));

    ----==== Loader signals ====----
    signal firmware_size            : std_logic_vector(RAM_ADDR_WIDTH + 2 downto 0) := (others => '0');
    signal loader_clk               : std_logic;
    signal loader_en_req            : std_logic;
    signal from_promless            : t_from_promless;
    signal loader_valid_pipe        : std_logic_vector(RAM_READ_LATENCY downto 0) := (others => '0');

    ------ Register signals begin (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    ------ Register signals end ----------------------------------------------
        
begin

    loader_clk <= to_promless_i.clk;
    loader_en_req <= to_promless_i.en;

    ----==== RAM instantiation ====----    

    i_gbtx_config_ram : xpm_memory_tdpram
        generic map(
            MEMORY_SIZE        => g_MAX_SIZE_BYTES * 8,
            MEMORY_PRIMITIVE   => g_MEMORY_PRIMITIVE,
            CLOCKING_MODE      => "common_clock",
            ECC_MODE           => "no_ecc",
            MEMORY_INIT_FILE   => "none",
            MEMORY_INIT_PARAM  => "0",
            USE_MEM_INIT       => 0,
            WAKEUP_TIME        => "disable_sleep",
            AUTO_SLEEP_TIME    => 0,
            MESSAGE_CONTROL    => 0,
            WRITE_DATA_WIDTH_A => 64,
            READ_DATA_WIDTH_A  => 64,
            BYTE_WRITE_WIDTH_A => 8,
            ADDR_WIDTH_A       => RAM_ADDR_WIDTH,
            READ_RESET_VALUE_A => "0",
            READ_LATENCY_A     => RAM_READ_LATENCY,
            WRITE_MODE_A       => "no_change",
            WRITE_DATA_WIDTH_B => 64,
            READ_DATA_WIDTH_B  => 64,
            BYTE_WRITE_WIDTH_B => 8,
            ADDR_WIDTH_B       => RAM_ADDR_WIDTH,
            READ_RESET_VALUE_B => "0",
            READ_LATENCY_B     => RAM_READ_LATENCY,
            WRITE_MODE_B       => "no_change"
        )
        port map(
            sleep          => '0',
            clka           => loader_clk,
            rsta           => '0',
            ena            => '1',
            regcea         => '1',
            wea            => rama_we,
            addra          => rama_addr,
            dina           => rama_din,
            injectsbiterra => '0',
            injectdbiterra => '0',
            douta          => rama_dout,
            sbiterra       => open,
            dbiterra       => open,
            clkb           => loader_clk,
            rstb           => '0',
            enb            => '1',
            regceb         => '1',
            web            => (others => '0'),
            addrb          => ramb_addr,
            dinb           => (others => '0'),
            injectsbiterrb => '0',
            injectdbiterrb => '0',
            doutb          => ramb_dout,
            sbiterrb       => open,
            dbiterrb       => open
        );

    ----==== BRAM reading / writing ====----    
    
    -- rama_din and rama_dout are connected to WRITE_DATA and READ_DATA registers
    -- whenever a write request to WRITE_DATA is done, WE is asserted and the write address is then incremented by 1
    -- same happens with the read requests
    process (loader_clk)
    begin
        if rising_edge(loader_clk) then
            if (reset_i = '1' or rama_reset_addr = '1') then
                rama_write_addr <= (others => '0');
                rama_read_addr <= (others => '0');
            else

                if (rama_write_req = '1') then
                    rama_addr <= rama_write_addr(RAM_ADDR_WIDTH downto 1);
                    -- select the upper or lower 32bit word based on the lowest address bit
                    if (rama_write_addr(0) = '0') then
                        rama_we <= x"0f";
                        rama_din <= x"00000000" & rama_write_data;
                    else
                        rama_we <= x"f0";
                        rama_din <= rama_write_data & x"00000000";
                    end if;
                elsif (rama_read_req = '1') then
                    rama_addr <= rama_read_addr(RAM_ADDR_WIDTH downto 1);
                    rama_we   <= (others => '0');
                    rama_din  <= (others => '0');
                else
                    rama_we   <= (others => '0');
                    rama_addr <= rama_addr;
                    rama_din  <= (others => '0');
                end if;
                
                -- increment the write address after WE has been asserted
                if (rama_we /= x"00") then
                    rama_write_addr <= std_logic_vector(unsigned(rama_write_addr) + 1);
                end if;

                -- increment the read address after read ready has been asserted
                if (rama_read_ready = '1') then
                    rama_read_addr <= std_logic_vector(unsigned(rama_read_addr) + 1);
                end if;
                
                -- delay the read ready signal
                rama_read_ready_pipe(0) <= rama_read_req;
                for i in 1 to RAM_READ_LATENCY loop
                    rama_read_ready_pipe(i) <= rama_read_ready_pipe(i - 1); 
                end loop;
                rama_read_ready <= rama_read_ready_pipe(RAM_READ_LATENCY);
                
                -- selct the upper or lower 32bit word based on the lowest bit of the read address
                if (rama_read_ready_pipe(RAM_READ_LATENCY) = '1') then
                    if (rama_read_addr(0) = '0') then
                        rama_read_data <= rama_dout(31 downto 0);
                    else
                        rama_read_data <= rama_dout(63 downto 32);
                    end if;
                end if;
                
            end if;
        end if;
    end process;

    ----==== Loader ====----    

    from_promless.first <= '0';
    from_promless.last <= '0';
    from_promless.error <= '0';

    process(loader_clk)
    begin
        if rising_edge(loader_clk) then
            if (reset_i = '1') then
                ramb_addr <= (others => '0');
                from_promless.ready <= '0';
                from_promless.valid <= '0';
                from_promless.data <= (others => '0');
                loader_valid_pipe <= (others => '0');
            else
                
                -- valid pipe
                for i in 1 to RAM_READ_LATENCY loop
                    loader_valid_pipe(i) <= loader_valid_pipe(i - 1); 
                end loop;
                from_promless.valid <= loader_valid_pipe(RAM_READ_LATENCY - 1);

                -- byte select pipe
                ramb_byte_sel_pipe(0) <= ramb_byte_sel;
                for i in 1 to RAM_READ_LATENCY loop
                    ramb_byte_sel_pipe(i) <= ramb_byte_sel_pipe(i - 1); 
                end loop;
                
                -- byte select
                case ramb_byte_sel_pipe(RAM_READ_LATENCY - 1) is
                    when "000" => from_promless.data <= ramb_dout(7 downto 0); 
                    when "001" => from_promless.data <= ramb_dout(15 downto 8); 
                    when "010" => from_promless.data <= ramb_dout(23 downto 16); 
                    when "011" => from_promless.data <= ramb_dout(31 downto 24); 
                    when "100" => from_promless.data <= ramb_dout(39 downto 32); 
                    when "101" => from_promless.data <= ramb_dout(47 downto 40); 
                    when "110" => from_promless.data <= ramb_dout(55 downto 48); 
                    when "111" => from_promless.data <= ramb_dout(63 downto 56); 
                end case;
                
                -- IDLE
                if (ramb_addr = std_logic_vector(to_unsigned(0, RAM_ADDR_WIDTH)) and ramb_byte_sel = "000") then
                    -- request
                    if (loader_en_req = '1') then
                        loader_valid_pipe(0) <= '1';
                        ramb_byte_sel <= std_logic_vector(unsigned(ramb_byte_sel) + 1);
                        ramb_addr <= ramb_addr;
                        from_promless.ready <= '0';
                    --idle
                    else
                        loader_valid_pipe(0) <= '0';
                        ramb_byte_sel <= "000";
                        ramb_addr <= (others => '0');
                        from_promless.ready <= '1';
                    end if;
                    
                -- DONE
                elsif (ramb_addr & ramb_byte_sel = firmware_size) then
                    loader_valid_pipe(0) <= '0';
                    ramb_addr <= (others => '0');
                    ramb_byte_sel <= (others => '0');
                    from_promless.ready <= '1';
                
                -- RUNNING
                else
                    loader_valid_pipe(0) <= '1';
                    from_promless.ready <= '0';
                    
                    if (ramb_byte_sel = "111") then
                        ramb_byte_sel <= "000";
                        ramb_addr <= std_logic_vector(unsigned(ramb_addr) + 1);
                    else
                        ramb_byte_sel <= std_logic_vector(unsigned(ramb_byte_sel) + 1);
                        ramb_addr <= ramb_addr;
                    end if;
                end if;
            end if;
        end if;
    end process;
        
    -- register the output
    process(loader_clk)
    begin
        if rising_edge(loader_clk) then
            from_promless_o <= from_promless;
        end if;
    end process;


    --===============================================================================================
    -- this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    --==== Registers end ============================================================================
    
end promless_arch;
